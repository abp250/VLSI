module add_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [15:0] A, B;
  output [16:0] Z;
  wire [15:0] A, B;
  wire [16:0] Z;
  wire n_51, n_56, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_134, n_135;
  nand g1 (n_51, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_56, A[1], B[1]);
  nand g10 (n_60, n_56, n_134, n_135);
  xor g11 (n_59, A[1], B[1]);
  nand g13 (n_61, A[2], B[2]);
  nand g14 (n_62, A[2], n_60);
  nand g15 (n_63, B[2], n_60);
  nand g16 (n_65, n_61, n_62, n_63);
  xor g17 (n_64, A[2], B[2]);
  xor g18 (Z[2], n_60, n_64);
  nand g19 (n_66, A[3], B[3]);
  nand g20 (n_67, A[3], n_65);
  nand g21 (n_68, B[3], n_65);
  nand g22 (n_70, n_66, n_67, n_68);
  xor g23 (n_69, A[3], B[3]);
  xor g24 (Z[3], n_65, n_69);
  nand g25 (n_71, A[4], B[4]);
  nand g26 (n_72, A[4], n_70);
  nand g27 (n_73, B[4], n_70);
  nand g28 (n_75, n_71, n_72, n_73);
  xor g29 (n_74, A[4], B[4]);
  xor g30 (Z[4], n_70, n_74);
  nand g31 (n_76, A[5], B[5]);
  nand g32 (n_77, A[5], n_75);
  nand g33 (n_78, B[5], n_75);
  nand g34 (n_80, n_76, n_77, n_78);
  xor g35 (n_79, A[5], B[5]);
  xor g36 (Z[5], n_75, n_79);
  nand g37 (n_81, A[6], B[6]);
  nand g38 (n_82, A[6], n_80);
  nand g39 (n_83, B[6], n_80);
  nand g40 (n_85, n_81, n_82, n_83);
  xor g41 (n_84, A[6], B[6]);
  xor g42 (Z[6], n_80, n_84);
  nand g43 (n_86, A[7], B[7]);
  nand g44 (n_87, A[7], n_85);
  nand g45 (n_88, B[7], n_85);
  nand g46 (n_90, n_86, n_87, n_88);
  xor g47 (n_89, A[7], B[7]);
  xor g48 (Z[7], n_85, n_89);
  nand g49 (n_91, A[8], B[8]);
  nand g50 (n_92, A[8], n_90);
  nand g51 (n_93, B[8], n_90);
  nand g52 (n_95, n_91, n_92, n_93);
  xor g53 (n_94, A[8], B[8]);
  xor g54 (Z[8], n_90, n_94);
  nand g55 (n_96, A[9], B[9]);
  nand g56 (n_97, A[9], n_95);
  nand g57 (n_98, B[9], n_95);
  nand g58 (n_100, n_96, n_97, n_98);
  xor g59 (n_99, A[9], B[9]);
  xor g60 (Z[9], n_95, n_99);
  nand g61 (n_101, A[10], B[10]);
  nand g62 (n_102, A[10], n_100);
  nand g63 (n_103, B[10], n_100);
  nand g64 (n_105, n_101, n_102, n_103);
  xor g65 (n_104, A[10], B[10]);
  xor g66 (Z[10], n_100, n_104);
  nand g67 (n_106, A[11], B[11]);
  nand g68 (n_107, A[11], n_105);
  nand g69 (n_108, B[11], n_105);
  nand g70 (n_110, n_106, n_107, n_108);
  xor g71 (n_109, A[11], B[11]);
  xor g72 (Z[11], n_105, n_109);
  nand g73 (n_111, A[12], B[12]);
  nand g74 (n_112, A[12], n_110);
  nand g75 (n_113, B[12], n_110);
  nand g76 (n_115, n_111, n_112, n_113);
  xor g77 (n_114, A[12], B[12]);
  xor g78 (Z[12], n_110, n_114);
  nand g79 (n_116, A[13], B[13]);
  nand g80 (n_117, A[13], n_115);
  nand g81 (n_118, B[13], n_115);
  nand g82 (n_120, n_116, n_117, n_118);
  xor g83 (n_119, A[13], B[13]);
  xor g84 (Z[13], n_115, n_119);
  nand g85 (n_121, A[14], B[14]);
  nand g86 (n_122, A[14], n_120);
  nand g87 (n_123, B[14], n_120);
  nand g88 (n_125, n_121, n_122, n_123);
  xor g89 (n_124, A[14], B[14]);
  xor g90 (Z[14], n_120, n_124);
  nand g91 (n_126, A[15], B[15]);
  nand g92 (n_127, A[15], n_125);
  nand g93 (n_128, B[15], n_125);
  nand g94 (Z[16], n_126, n_127, n_128);
  xor g95 (n_129, A[15], B[15]);
  xor g96 (Z[15], n_125, n_129);
  or g98 (n_134, wc, n_51);
  not gc (wc, A[1]);
  or g99 (n_135, wc0, n_51);
  not gc0 (wc0, B[1]);
  xnor g100 (Z[1], n_51, n_59);
endmodule

module add_unsigned_GENERIC(A, B, Z);
  input [15:0] A, B;
  output [16:0] Z;
  wire [15:0] A, B;
  wire [16:0] Z;
  add_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_162_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [16:0] A, B;
  output [16:0] Z;
  wire [16:0] A, B;
  wire [16:0] Z;
  wire n_53, n_58, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_136, n_142, n_143;
  nand g1 (n_53, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_58, A[1], B[1]);
  nand g10 (n_62, n_58, n_142, n_143);
  xor g11 (n_61, A[1], B[1]);
  nand g13 (n_63, A[2], B[2]);
  nand g14 (n_64, A[2], n_62);
  nand g15 (n_65, B[2], n_62);
  nand g16 (n_67, n_63, n_64, n_65);
  xor g17 (n_66, A[2], B[2]);
  xor g18 (Z[2], n_62, n_66);
  nand g19 (n_68, A[3], B[3]);
  nand g20 (n_69, A[3], n_67);
  nand g21 (n_70, B[3], n_67);
  nand g22 (n_72, n_68, n_69, n_70);
  xor g23 (n_71, A[3], B[3]);
  xor g24 (Z[3], n_67, n_71);
  nand g25 (n_73, A[4], B[4]);
  nand g26 (n_74, A[4], n_72);
  nand g27 (n_75, B[4], n_72);
  nand g28 (n_77, n_73, n_74, n_75);
  xor g29 (n_76, A[4], B[4]);
  xor g30 (Z[4], n_72, n_76);
  nand g31 (n_78, A[5], B[5]);
  nand g32 (n_79, A[5], n_77);
  nand g33 (n_80, B[5], n_77);
  nand g34 (n_82, n_78, n_79, n_80);
  xor g35 (n_81, A[5], B[5]);
  xor g36 (Z[5], n_77, n_81);
  nand g37 (n_83, A[6], B[6]);
  nand g38 (n_84, A[6], n_82);
  nand g39 (n_85, B[6], n_82);
  nand g40 (n_87, n_83, n_84, n_85);
  xor g41 (n_86, A[6], B[6]);
  xor g42 (Z[6], n_82, n_86);
  nand g43 (n_88, A[7], B[7]);
  nand g44 (n_89, A[7], n_87);
  nand g45 (n_90, B[7], n_87);
  nand g46 (n_92, n_88, n_89, n_90);
  xor g47 (n_91, A[7], B[7]);
  xor g48 (Z[7], n_87, n_91);
  nand g49 (n_93, A[8], B[8]);
  nand g50 (n_94, A[8], n_92);
  nand g51 (n_95, B[8], n_92);
  nand g52 (n_97, n_93, n_94, n_95);
  xor g53 (n_96, A[8], B[8]);
  xor g54 (Z[8], n_92, n_96);
  nand g55 (n_98, A[9], B[9]);
  nand g56 (n_99, A[9], n_97);
  nand g57 (n_100, B[9], n_97);
  nand g58 (n_102, n_98, n_99, n_100);
  xor g59 (n_101, A[9], B[9]);
  xor g60 (Z[9], n_97, n_101);
  nand g61 (n_103, A[10], B[10]);
  nand g62 (n_104, A[10], n_102);
  nand g63 (n_105, B[10], n_102);
  nand g64 (n_107, n_103, n_104, n_105);
  xor g65 (n_106, A[10], B[10]);
  xor g66 (Z[10], n_102, n_106);
  nand g67 (n_108, A[11], B[11]);
  nand g68 (n_109, A[11], n_107);
  nand g69 (n_110, B[11], n_107);
  nand g70 (n_112, n_108, n_109, n_110);
  xor g71 (n_111, A[11], B[11]);
  xor g72 (Z[11], n_107, n_111);
  nand g73 (n_113, A[12], B[12]);
  nand g74 (n_114, A[12], n_112);
  nand g75 (n_115, B[12], n_112);
  nand g76 (n_117, n_113, n_114, n_115);
  xor g77 (n_116, A[12], B[12]);
  xor g78 (Z[12], n_112, n_116);
  nand g79 (n_118, A[13], B[13]);
  nand g80 (n_119, A[13], n_117);
  nand g81 (n_120, B[13], n_117);
  nand g82 (n_122, n_118, n_119, n_120);
  xor g83 (n_121, A[13], B[13]);
  xor g84 (Z[13], n_117, n_121);
  nand g85 (n_123, A[14], B[14]);
  nand g86 (n_124, A[14], n_122);
  nand g87 (n_125, B[14], n_122);
  nand g88 (n_127, n_123, n_124, n_125);
  xor g89 (n_126, A[14], B[14]);
  xor g90 (Z[14], n_122, n_126);
  nand g91 (n_128, A[15], B[15]);
  nand g92 (n_129, A[15], n_127);
  nand g93 (n_130, B[15], n_127);
  nand g94 (n_132, n_128, n_129, n_130);
  xor g95 (n_131, A[15], B[15]);
  xor g96 (Z[15], n_127, n_131);
  xor g101 (n_136, A[16], B[16]);
  xor g102 (Z[16], n_132, n_136);
  or g104 (n_142, wc, n_53);
  not gc (wc, A[1]);
  or g105 (n_143, wc0, n_53);
  not gc0 (wc0, B[1]);
  xnor g106 (Z[1], n_53, n_61);
endmodule

module add_unsigned_162_GENERIC(A, B, Z);
  input [16:0] A, B;
  output [16:0] Z;
  wire [16:0] A, B;
  wire [16:0] Z;
  add_unsigned_162_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module mult_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $unsigned(A) * $unsigned(B);"
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_325;
  wire n_328, n_330, n_333, n_335, n_336, n_338, n_340, n_341;
  wire n_343, n_345, n_346, n_348, n_350, n_351, n_353, n_355;
  wire n_356, n_358, n_360, n_361, n_363, n_365, n_366, n_368;
  wire n_370, n_371, n_373, n_375, n_376, n_378, n_380, n_381;
  wire n_383, n_385, n_386, n_388, n_390, n_391, n_393, n_417;
  wire n_419, n_420, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445;
  and g1 (Z[0], A[0], B[0]);
  and g2 (n_46, A[1], B[0]);
  and g3 (n_63, A[2], B[0]);
  and g4 (n_67, A[3], B[0]);
  and g5 (n_72, A[4], B[0]);
  and g6 (n_80, A[5], B[0]);
  and g7 (n_90, A[6], B[0]);
  and g8 (n_103, A[7], B[0]);
  and g9 (n_61, A[0], B[1]);
  and g10 (n_45, A[1], B[1]);
  and g11 (n_68, A[2], B[1]);
  and g12 (n_73, A[3], B[1]);
  and g13 (n_64, A[4], B[1]);
  and g14 (n_91, A[5], B[1]);
  and g15 (n_104, A[6], B[1]);
  and g16 (n_120, A[7], B[1]);
  and g17 (n_66, A[0], B[2]);
  and g18 (n_70, A[1], B[2]);
  and g19 (n_76, A[2], B[2]);
  and g20 (n_83, A[3], B[2]);
  and g21 (n_94, A[4], B[2]);
  and g22 (n_108, A[5], B[2]);
  and g23 (n_121, A[6], B[2]);
  and g24 (n_137, A[7], B[2]);
  and g25 (n_69, A[0], B[3]);
  and g26 (n_74, A[1], B[3]);
  and g27 (n_81, A[2], B[3]);
  and g28 (n_92, A[3], B[3]);
  and g29 (n_105, A[4], B[3]);
  and g30 (n_124, A[5], B[3]);
  and g31 (n_138, A[6], B[3]);
  and g32 (n_152, A[7], B[3]);
  and g33 (n_75, A[0], B[4]);
  and g34 (n_82, A[1], B[4]);
  and g35 (n_93, A[2], B[4]);
  and g36 (n_107, A[3], B[4]);
  and g37 (n_122, A[4], B[4]);
  and g38 (n_141, A[5], B[4]);
  and g39 (n_153, A[6], B[4]);
  and g40 (n_164, A[7], B[4]);
  and g41 (n_84, A[0], B[5]);
  and g42 (n_65, A[1], B[5]);
  and g43 (n_109, A[2], B[5]);
  and g44 (n_123, A[3], B[5]);
  and g45 (n_139, A[4], B[5]);
  and g46 (n_156, A[5], B[5]);
  and g47 (n_165, A[6], B[5]);
  and g48 (n_173, A[7], B[5]);
  and g49 (n_95, A[0], B[6]);
  and g50 (n_110, A[1], B[6]);
  and g51 (n_125, A[2], B[6]);
  and g52 (n_140, A[3], B[6]);
  and g53 (n_154, A[4], B[6]);
  and g54 (n_167, A[5], B[6]);
  and g55 (n_174, A[6], B[6]);
  and g56 (n_179, A[7], B[6]);
  and g57 (n_106, A[0], B[7]);
  and g58 (n_126, A[1], B[7]);
  and g59 (n_142, A[2], B[7]);
  and g60 (n_155, A[3], B[7]);
  and g61 (n_166, A[4], B[7]);
  and g62 (n_175, A[5], B[7]);
  and g63 (n_180, A[6], B[7]);
  and g64 (n_33, A[7], B[7]);
  xor g107 (n_60, n_63, n_66);
  and g108 (n_44, n_63, n_66);
  xor g109 (n_71, n_67, n_68);
  and g110 (n_78, n_67, n_68);
  xor g111 (n_182, n_69, n_70);
  xor g112 (n_59, n_182, n_71);
  nand g113 (n_183, n_69, n_70);
  nand g114 (n_184, n_71, n_70);
  nand g115 (n_185, n_69, n_71);
  nand g116 (n_43, n_183, n_184, n_185);
  xor g117 (n_77, n_72, n_73);
  and g118 (n_86, n_72, n_73);
  xor g119 (n_186, n_74, n_75);
  xor g120 (n_79, n_186, n_76);
  nand g121 (n_187, n_74, n_75);
  nand g122 (n_188, n_76, n_75);
  nand g123 (n_189, n_74, n_76);
  nand g124 (n_87, n_187, n_188, n_189);
  xor g125 (n_190, n_77, n_78);
  xor g126 (n_58, n_190, n_79);
  nand g127 (n_191, n_77, n_78);
  nand g128 (n_192, n_79, n_78);
  nand g129 (n_193, n_77, n_79);
  nand g130 (n_42, n_191, n_192, n_193);
  xor g131 (n_85, n_80, n_64);
  and g132 (n_96, n_80, n_64);
  xor g133 (n_194, n_81, n_82);
  xor g134 (n_88, n_194, n_83);
  nand g135 (n_195, n_81, n_82);
  nand g136 (n_196, n_83, n_82);
  nand g137 (n_197, n_81, n_83);
  nand g138 (n_98, n_195, n_196, n_197);
  xor g139 (n_198, n_84, n_85);
  xor g140 (n_89, n_198, n_86);
  nand g141 (n_199, n_84, n_85);
  nand g142 (n_200, n_86, n_85);
  nand g143 (n_201, n_84, n_86);
  nand g144 (n_100, n_199, n_200, n_201);
  xor g145 (n_202, n_87, n_88);
  xor g146 (n_57, n_202, n_89);
  nand g147 (n_203, n_87, n_88);
  nand g148 (n_204, n_89, n_88);
  nand g149 (n_205, n_87, n_89);
  nand g150 (n_41, n_203, n_204, n_205);
  xor g151 (n_97, n_90, n_91);
  and g152 (n_111, n_90, n_91);
  xor g153 (n_206, n_92, n_93);
  xor g154 (n_99, n_206, n_94);
  nand g155 (n_207, n_92, n_93);
  nand g156 (n_208, n_94, n_93);
  nand g157 (n_209, n_92, n_94);
  nand g158 (n_113, n_207, n_208, n_209);
  xor g159 (n_210, n_65, n_95);
  xor g160 (n_101, n_210, n_96);
  nand g161 (n_211, n_65, n_95);
  nand g162 (n_212, n_96, n_95);
  nand g163 (n_213, n_65, n_96);
  nand g164 (n_116, n_211, n_212, n_213);
  xor g165 (n_214, n_97, n_98);
  xor g166 (n_102, n_214, n_99);
  nand g167 (n_215, n_97, n_98);
  nand g168 (n_216, n_99, n_98);
  nand g169 (n_217, n_97, n_99);
  nand g170 (n_118, n_215, n_216, n_217);
  xor g171 (n_218, n_100, n_101);
  xor g172 (n_56, n_218, n_102);
  nand g173 (n_219, n_100, n_101);
  nand g174 (n_220, n_102, n_101);
  nand g175 (n_221, n_100, n_102);
  nand g176 (n_40, n_219, n_220, n_221);
  xor g177 (n_112, n_103, n_104);
  and g178 (n_128, n_103, n_104);
  xor g179 (n_222, n_105, n_106);
  xor g180 (n_115, n_222, n_107);
  nand g181 (n_223, n_105, n_106);
  nand g182 (n_224, n_107, n_106);
  nand g183 (n_225, n_105, n_107);
  nand g184 (n_129, n_223, n_224, n_225);
  xor g185 (n_226, n_108, n_109);
  xor g186 (n_114, n_226, n_110);
  nand g187 (n_227, n_108, n_109);
  nand g188 (n_228, n_110, n_109);
  nand g189 (n_229, n_108, n_110);
  nand g190 (n_130, n_227, n_228, n_229);
  xor g191 (n_230, n_111, n_112);
  xor g192 (n_117, n_230, n_113);
  nand g193 (n_231, n_111, n_112);
  nand g194 (n_232, n_113, n_112);
  nand g195 (n_233, n_111, n_113);
  nand g196 (n_133, n_231, n_232, n_233);
  xor g197 (n_234, n_114, n_115);
  xor g198 (n_119, n_234, n_116);
  nand g199 (n_235, n_114, n_115);
  nand g200 (n_236, n_116, n_115);
  nand g201 (n_237, n_114, n_116);
  nand g202 (n_135, n_235, n_236, n_237);
  xor g203 (n_238, n_117, n_118);
  xor g204 (n_55, n_238, n_119);
  nand g205 (n_239, n_117, n_118);
  nand g206 (n_240, n_119, n_118);
  nand g207 (n_241, n_117, n_119);
  nand g208 (n_39, n_239, n_240, n_241);
  xor g209 (n_127, n_120, n_121);
  and g210 (n_143, n_120, n_121);
  xor g211 (n_242, n_122, n_123);
  xor g212 (n_131, n_242, n_124);
  nand g213 (n_243, n_122, n_123);
  nand g214 (n_244, n_124, n_123);
  nand g215 (n_245, n_122, n_124);
  nand g216 (n_144, n_243, n_244, n_245);
  xor g217 (n_246, n_125, n_126);
  xor g218 (n_132, n_246, n_127);
  nand g219 (n_247, n_125, n_126);
  nand g220 (n_248, n_127, n_126);
  nand g221 (n_249, n_125, n_127);
  nand g222 (n_147, n_247, n_248, n_249);
  xor g223 (n_250, n_128, n_129);
  xor g224 (n_134, n_250, n_130);
  nand g225 (n_251, n_128, n_129);
  nand g226 (n_252, n_130, n_129);
  nand g227 (n_253, n_128, n_130);
  nand g228 (n_148, n_251, n_252, n_253);
  xor g229 (n_254, n_131, n_132);
  xor g230 (n_136, n_254, n_133);
  nand g231 (n_255, n_131, n_132);
  nand g232 (n_256, n_133, n_132);
  nand g233 (n_257, n_131, n_133);
  nand g234 (n_151, n_255, n_256, n_257);
  xor g235 (n_258, n_134, n_135);
  xor g236 (n_54, n_258, n_136);
  nand g237 (n_259, n_134, n_135);
  nand g238 (n_260, n_136, n_135);
  nand g239 (n_261, n_134, n_136);
  nand g240 (n_38, n_259, n_260, n_261);
  xor g241 (n_262, n_137, n_138);
  xor g242 (n_146, n_262, n_139);
  nand g243 (n_263, n_137, n_138);
  nand g244 (n_264, n_139, n_138);
  nand g245 (n_265, n_137, n_139);
  nand g246 (n_158, n_263, n_264, n_265);
  xor g247 (n_266, n_140, n_141);
  xor g248 (n_145, n_266, n_142);
  nand g249 (n_267, n_140, n_141);
  nand g250 (n_268, n_142, n_141);
  nand g251 (n_269, n_140, n_142);
  nand g252 (n_157, n_267, n_268, n_269);
  xor g253 (n_270, n_143, n_144);
  xor g254 (n_149, n_270, n_145);
  nand g255 (n_271, n_143, n_144);
  nand g256 (n_272, n_145, n_144);
  nand g257 (n_273, n_143, n_145);
  nand g258 (n_161, n_271, n_272, n_273);
  xor g259 (n_274, n_146, n_147);
  xor g260 (n_150, n_274, n_148);
  nand g261 (n_275, n_146, n_147);
  nand g262 (n_276, n_148, n_147);
  nand g263 (n_277, n_146, n_148);
  nand g264 (n_163, n_275, n_276, n_277);
  xor g265 (n_278, n_149, n_150);
  xor g266 (n_53, n_278, n_151);
  nand g267 (n_279, n_149, n_150);
  nand g268 (n_280, n_151, n_150);
  nand g269 (n_281, n_149, n_151);
  nand g270 (n_37, n_279, n_280, n_281);
  xor g271 (n_282, n_152, n_153);
  xor g272 (n_159, n_282, n_154);
  nand g273 (n_283, n_152, n_153);
  nand g274 (n_284, n_154, n_153);
  nand g275 (n_285, n_152, n_154);
  nand g276 (n_168, n_283, n_284, n_285);
  xor g277 (n_286, n_155, n_156);
  xor g278 (n_160, n_286, n_157);
  nand g279 (n_287, n_155, n_156);
  nand g280 (n_288, n_157, n_156);
  nand g281 (n_289, n_155, n_157);
  nand g282 (n_170, n_287, n_288, n_289);
  xor g283 (n_290, n_158, n_159);
  xor g284 (n_162, n_290, n_160);
  nand g285 (n_291, n_158, n_159);
  nand g286 (n_292, n_160, n_159);
  nand g287 (n_293, n_158, n_160);
  nand g288 (n_172, n_291, n_292, n_293);
  xor g289 (n_294, n_161, n_162);
  xor g290 (n_52, n_294, n_163);
  nand g291 (n_295, n_161, n_162);
  nand g292 (n_296, n_163, n_162);
  nand g293 (n_297, n_161, n_163);
  nand g294 (n_36, n_295, n_296, n_297);
  xor g295 (n_298, n_164, n_165);
  xor g296 (n_169, n_298, n_166);
  nand g297 (n_299, n_164, n_165);
  nand g298 (n_300, n_166, n_165);
  nand g299 (n_301, n_164, n_166);
  nand g300 (n_176, n_299, n_300, n_301);
  xor g301 (n_302, n_167, n_168);
  xor g302 (n_171, n_302, n_169);
  nand g303 (n_303, n_167, n_168);
  nand g304 (n_304, n_169, n_168);
  nand g305 (n_305, n_167, n_169);
  nand g306 (n_178, n_303, n_304, n_305);
  xor g307 (n_306, n_170, n_171);
  xor g308 (n_51, n_306, n_172);
  nand g309 (n_307, n_170, n_171);
  nand g310 (n_308, n_172, n_171);
  nand g311 (n_309, n_170, n_172);
  nand g312 (n_50, n_307, n_308, n_309);
  xor g313 (n_310, n_173, n_174);
  xor g314 (n_177, n_310, n_175);
  nand g315 (n_311, n_173, n_174);
  nand g316 (n_312, n_175, n_174);
  nand g317 (n_313, n_173, n_175);
  nand g318 (n_181, n_311, n_312, n_313);
  xor g319 (n_314, n_176, n_177);
  xor g320 (n_35, n_314, n_178);
  nand g321 (n_315, n_176, n_177);
  nand g322 (n_316, n_178, n_177);
  nand g323 (n_317, n_176, n_178);
  nand g324 (n_49, n_315, n_316, n_317);
  xor g325 (n_318, n_179, n_180);
  xor g326 (n_34, n_318, n_181);
  nand g327 (n_319, n_179, n_180);
  nand g328 (n_320, n_181, n_180);
  nand g329 (n_321, n_179, n_181);
  nand g330 (n_48, n_319, n_320, n_321);
  nor g336 (n_325, n_46, n_61);
  nand g337 (n_328, n_46, n_61);
  nor g338 (n_330, n_45, n_60);
  nand g339 (n_333, n_45, n_60);
  nor g340 (n_335, n_44, n_59);
  nand g341 (n_338, n_44, n_59);
  nor g342 (n_340, n_43, n_58);
  nand g343 (n_343, n_43, n_58);
  nor g344 (n_345, n_42, n_57);
  nand g345 (n_348, n_42, n_57);
  nor g346 (n_350, n_41, n_56);
  nand g347 (n_353, n_41, n_56);
  nor g348 (n_355, n_40, n_55);
  nand g349 (n_358, n_40, n_55);
  nor g350 (n_360, n_39, n_54);
  nand g351 (n_363, n_39, n_54);
  nor g352 (n_365, n_38, n_53);
  nand g353 (n_368, n_38, n_53);
  nor g354 (n_370, n_37, n_52);
  nand g355 (n_373, n_37, n_52);
  nor g356 (n_375, n_36, n_51);
  nand g357 (n_378, n_36, n_51);
  nor g358 (n_380, n_35, n_50);
  nand g359 (n_383, n_35, n_50);
  nor g360 (n_385, n_34, n_49);
  nand g361 (n_388, n_34, n_49);
  nor g362 (n_390, n_33, n_48);
  nand g363 (n_393, n_33, n_48);
  nand g371 (n_336, n_333, n_420);
  nand g374 (n_341, n_338, n_424);
  nand g377 (n_346, n_343, n_428);
  nand g380 (n_351, n_348, n_434);
  nand g383 (n_356, n_353, n_437);
  nand g386 (n_361, n_358, n_438);
  nand g389 (n_366, n_363, n_439);
  nand g392 (n_371, n_368, n_440);
  nand g65 (n_376, n_373, n_441);
  nand g68 (n_381, n_378, n_442);
  nand g71 (n_386, n_383, n_443);
  nand g74 (n_391, n_388, n_444);
  nand g77 (Z[15], n_393, n_445);
  xnor g86 (Z[3], n_336, n_422);
  xnor g88 (Z[4], n_341, n_423);
  xnor g90 (Z[5], n_346, n_425);
  xnor g92 (Z[6], n_351, n_427);
  xnor g94 (Z[7], n_356, n_429);
  xnor g96 (Z[8], n_361, n_431);
  xnor g98 (Z[9], n_366, n_432);
  xnor g100 (Z[10], n_371, n_435);
  xnor g102 (Z[11], n_376, n_436);
  xnor g104 (Z[12], n_381, n_433);
  xnor g106 (Z[13], n_386, n_430);
  xnor g396 (Z[14], n_391, n_426);
  or g400 (n_417, wc, n_325);
  not gc (wc, n_328);
  not g402 (Z[1], n_417);
  or g403 (n_419, wc0, n_330);
  not gc0 (wc0, n_333);
  or g404 (n_420, n_328, n_330);
  xor g405 (Z[2], n_328, n_419);
  or g406 (n_422, wc1, n_335);
  not gc1 (wc1, n_338);
  or g407 (n_423, wc2, n_340);
  not gc2 (wc2, n_343);
  or g408 (n_424, wc3, n_335);
  not gc3 (wc3, n_336);
  or g409 (n_425, wc4, n_345);
  not gc4 (wc4, n_348);
  or g410 (n_426, wc5, n_390);
  not gc5 (wc5, n_393);
  or g411 (n_427, wc6, n_350);
  not gc6 (wc6, n_353);
  or g412 (n_428, wc7, n_340);
  not gc7 (wc7, n_341);
  or g413 (n_429, wc8, n_355);
  not gc8 (wc8, n_358);
  or g414 (n_430, wc9, n_385);
  not gc9 (wc9, n_388);
  or g415 (n_431, wc10, n_360);
  not gc10 (wc10, n_363);
  or g416 (n_432, wc11, n_365);
  not gc11 (wc11, n_368);
  or g417 (n_433, wc12, n_380);
  not gc12 (wc12, n_383);
  or g418 (n_434, wc13, n_345);
  not gc13 (wc13, n_346);
  or g419 (n_435, wc14, n_370);
  not gc14 (wc14, n_373);
  or g420 (n_436, wc15, n_375);
  not gc15 (wc15, n_378);
  or g421 (n_437, wc16, n_350);
  not gc16 (wc16, n_351);
  or g422 (n_438, wc17, n_355);
  not gc17 (wc17, n_356);
  or g423 (n_439, wc18, n_360);
  not gc18 (wc18, n_361);
  or g424 (n_440, wc19, n_365);
  not gc19 (wc19, n_366);
  or g425 (n_441, wc20, n_370);
  not gc20 (wc20, n_371);
  or g426 (n_442, wc21, n_375);
  not gc21 (wc21, n_376);
  or g427 (n_443, wc22, n_380);
  not gc22 (wc22, n_381);
  or g428 (n_444, wc23, n_385);
  not gc23 (wc23, n_386);
  or g429 (n_445, wc24, n_390);
  not gc24 (wc24, n_391);
endmodule

module mult_unsigned_GENERIC(A, B, Z);
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  mult_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module mult_unsigned_120_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $unsigned(A) * $unsigned(B);"
  input [15:0] A, B;
  output [16:0] Z;
  wire [15:0] A, B;
  wire [16:0] Z;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_84, n_87, n_88, n_89, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_138, n_139, n_145, n_147, n_148, n_149, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_196, n_198, n_199, n_200, n_202, n_203, n_204, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_245, n_247, n_248, n_249, n_251;
  wire n_252, n_253, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_288, n_290, n_291, n_292, n_294, n_295, n_296, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316;
  wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_325;
  wire n_327, n_328, n_329, n_331, n_332, n_333, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_356, n_358, n_359, n_360, n_362, n_363, n_364, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_381, n_383, n_384, n_385, n_387;
  wire n_388, n_389, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_400, n_402, n_403, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584;
  wire n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592;
  wire n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672;
  wire n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696;
  wire n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704;
  wire n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_745, n_749, n_753;
  wire n_757, n_761, n_765, n_774, n_777, n_779, n_782, n_784;
  wire n_785, n_787, n_789, n_790, n_792, n_794, n_795, n_797;
  wire n_799, n_800, n_802, n_804, n_805, n_807, n_809, n_810;
  wire n_812, n_814, n_815, n_817, n_819, n_820, n_822, n_824;
  wire n_825, n_827, n_829, n_830, n_832, n_834, n_835, n_837;
  wire n_839, n_840, n_842, n_844, n_845, n_847, n_850, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_882, n_883;
  wire n_885, n_886, n_888, n_889, n_890, n_891, n_892, n_893;
  wire n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901;
  wire n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909;
  wire n_910, n_911, n_912, n_913, n_914, n_915;
  xor g2 (n_87, B[1], B[0]);
  xor g8 (n_88, B[1], A[0]);
  and g12 (Z[0], A[0], B[0]);
  xor g13 (n_93, B[1], A[1]);
  nand g14 (n_94, n_93, B[0]);
  nand g15 (n_95, n_88, n_89);
  nand g16 (n_82, n_94, n_95);
  xor g17 (n_96, B[1], A[2]);
  nand g18 (n_97, n_96, B[0]);
  nand g19 (n_98, n_93, n_89);
  nand g20 (n_81, n_97, n_98);
  xor g21 (n_99, B[1], A[3]);
  nand g22 (n_100, n_99, B[0]);
  nand g23 (n_101, n_96, n_89);
  nand g24 (n_413, n_100, n_101);
  xor g25 (n_102, B[1], A[4]);
  nand g26 (n_103, n_102, B[0]);
  nand g27 (n_104, n_99, n_89);
  nand g28 (n_414, n_103, n_104);
  xor g29 (n_105, B[1], A[5]);
  nand g30 (n_106, n_105, B[0]);
  nand g31 (n_107, n_102, n_89);
  nand g32 (n_419, n_106, n_107);
  xor g33 (n_108, B[1], A[6]);
  nand g34 (n_109, n_108, B[0]);
  nand g35 (n_110, n_105, n_89);
  nand g36 (n_425, n_109, n_110);
  xor g37 (n_111, B[1], A[7]);
  nand g38 (n_112, n_111, B[0]);
  nand g39 (n_113, n_108, n_89);
  nand g40 (n_430, n_112, n_113);
  xor g41 (n_114, B[1], A[8]);
  nand g42 (n_115, n_114, B[0]);
  nand g43 (n_116, n_111, n_89);
  nand g44 (n_440, n_115, n_116);
  xor g45 (n_117, B[1], A[9]);
  nand g46 (n_118, n_117, B[0]);
  nand g47 (n_119, n_114, n_89);
  nand g48 (n_450, n_118, n_119);
  xor g49 (n_120, B[1], A[10]);
  nand g50 (n_121, n_120, B[0]);
  nand g51 (n_122, n_117, n_89);
  nand g52 (n_460, n_121, n_122);
  xor g53 (n_123, B[1], A[11]);
  nand g54 (n_124, n_123, B[0]);
  nand g55 (n_125, n_120, n_89);
  nand g56 (n_472, n_124, n_125);
  xor g57 (n_126, B[1], A[12]);
  nand g58 (n_127, n_126, B[0]);
  nand g59 (n_128, n_123, n_89);
  nand g60 (n_486, n_127, n_128);
  xor g61 (n_129, B[1], A[13]);
  nand g62 (n_130, n_129, B[0]);
  nand g63 (n_131, n_126, n_89);
  nand g64 (n_503, n_130, n_131);
  xor g65 (n_84, B[1], A[14]);
  nand g66 (n_132, n_84, B[0]);
  nand g67 (n_133, n_129, n_89);
  nand g68 (n_519, n_132, n_133);
  xor g69 (n_134, B[1], A[15]);
  nand g70 (n_135, n_134, B[0]);
  nand g71 (n_136, n_84, n_89);
  nand g72 (n_537, n_135, n_136);
  nand g74 (n_138, B[1], B[0]);
  nand g75 (n_139, n_134, n_89);
  nand g76 (n_557, n_138, n_139);
  xor g81 (n_145, B[2], B[1]);
  xor g82 (n_147, B[3], B[2]);
  nor g86 (n_198, B[1], B[2]);
  nand g87 (n_196, B[1], B[2]);
  xor g88 (n_148, B[3], A[0]);
  and g92 (n_64, A[0], n_145);
  xor g93 (n_153, B[3], A[1]);
  nand g94 (n_154, n_153, n_145);
  nand g95 (n_155, n_148, n_149);
  nand g96 (n_63, n_154, n_155);
  xor g97 (n_156, B[3], A[2]);
  nand g98 (n_157, n_156, n_145);
  nand g99 (n_158, n_153, n_149);
  nand g100 (n_415, n_157, n_158);
  xor g101 (n_159, B[3], A[3]);
  nand g102 (n_160, n_159, n_145);
  nand g103 (n_161, n_156, n_149);
  nand g104 (n_417, n_160, n_161);
  xor g105 (n_162, B[3], A[4]);
  nand g106 (n_163, n_162, n_145);
  nand g107 (n_164, n_159, n_149);
  nand g108 (n_422, n_163, n_164);
  xor g109 (n_165, B[3], A[5]);
  nand g110 (n_166, n_165, n_145);
  nand g111 (n_167, n_162, n_149);
  nand g112 (n_429, n_166, n_167);
  xor g113 (n_168, B[3], A[6]);
  nand g114 (n_169, n_168, n_145);
  nand g115 (n_170, n_165, n_149);
  nand g116 (n_436, n_169, n_170);
  xor g117 (n_171, B[3], A[7]);
  nand g118 (n_172, n_171, n_145);
  nand g119 (n_173, n_168, n_149);
  nand g120 (n_445, n_172, n_173);
  xor g121 (n_174, B[3], A[8]);
  nand g122 (n_175, n_174, n_145);
  nand g123 (n_176, n_171, n_149);
  nand g124 (n_458, n_175, n_176);
  xor g125 (n_177, B[3], A[9]);
  nand g126 (n_178, n_177, n_145);
  nand g127 (n_179, n_174, n_149);
  nand g128 (n_471, n_178, n_179);
  xor g129 (n_180, B[3], A[10]);
  nand g130 (n_181, n_180, n_145);
  nand g131 (n_182, n_177, n_149);
  nand g132 (n_484, n_181, n_182);
  xor g133 (n_183, B[3], A[11]);
  nand g134 (n_184, n_183, n_145);
  nand g135 (n_185, n_180, n_149);
  nand g136 (n_501, n_184, n_185);
  xor g137 (n_186, B[3], A[12]);
  nand g138 (n_187, n_186, n_145);
  nand g139 (n_188, n_183, n_149);
  nand g140 (n_518, n_187, n_188);
  xor g141 (n_189, B[3], A[13]);
  nand g142 (n_190, n_189, n_145);
  nand g143 (n_191, n_186, n_149);
  nand g144 (n_536, n_190, n_191);
  xor g145 (n_192, B[3], A[14]);
  nand g146 (n_193, n_192, n_145);
  nand g147 (n_194, n_189, n_149);
  nand g148 (n_556, n_193, n_194);
  or g151 (n_199, n_873, n_198);
  and g152 (n_412, B[3], n_199);
  xor g153 (n_200, B[4], B[3]);
  xor g154 (n_202, B[5], B[4]);
  nor g158 (n_247, B[3], B[4]);
  nand g159 (n_245, B[3], B[4]);
  xor g160 (n_203, B[5], A[0]);
  and g164 (n_416, A[0], n_200);
  xor g165 (n_208, B[5], A[1]);
  nand g166 (n_209, n_208, n_200);
  nand g167 (n_210, n_203, n_204);
  nand g168 (n_421, n_209, n_210);
  xor g169 (n_211, B[5], A[2]);
  nand g170 (n_212, n_211, n_200);
  nand g171 (n_213, n_208, n_204);
  nand g172 (n_426, n_212, n_213);
  xor g173 (n_214, B[5], A[3]);
  nand g174 (n_215, n_214, n_200);
  nand g175 (n_216, n_211, n_204);
  nand g176 (n_431, n_215, n_216);
  xor g177 (n_217, B[5], A[4]);
  nand g178 (n_218, n_217, n_200);
  nand g179 (n_219, n_214, n_204);
  nand g180 (n_438, n_218, n_219);
  xor g181 (n_220, B[5], A[5]);
  nand g182 (n_221, n_220, n_200);
  nand g183 (n_222, n_217, n_204);
  nand g184 (n_446, n_221, n_222);
  xor g185 (n_223, B[5], A[6]);
  nand g186 (n_224, n_223, n_200);
  nand g187 (n_225, n_220, n_204);
  nand g188 (n_456, n_224, n_225);
  xor g189 (n_226, B[5], A[7]);
  nand g190 (n_227, n_226, n_200);
  nand g191 (n_228, n_223, n_204);
  nand g192 (n_468, n_227, n_228);
  xor g193 (n_229, B[5], A[8]);
  nand g194 (n_230, n_229, n_200);
  nand g195 (n_231, n_226, n_204);
  nand g196 (n_482, n_230, n_231);
  xor g197 (n_232, B[5], A[9]);
  nand g198 (n_233, n_232, n_200);
  nand g199 (n_234, n_229, n_204);
  nand g200 (n_498, n_233, n_234);
  xor g201 (n_235, B[5], A[10]);
  nand g202 (n_236, n_235, n_200);
  nand g203 (n_237, n_232, n_204);
  nand g204 (n_515, n_236, n_237);
  xor g205 (n_238, B[5], A[11]);
  nand g206 (n_239, n_238, n_200);
  nand g207 (n_240, n_235, n_204);
  nand g208 (n_533, n_239, n_240);
  xor g209 (n_241, B[5], A[12]);
  nand g210 (n_242, n_241, n_200);
  nand g211 (n_243, n_238, n_204);
  nand g212 (n_553, n_242, n_243);
  or g215 (n_248, n_874, n_247);
  and g216 (n_418, B[5], n_248);
  xor g217 (n_249, B[6], B[5]);
  xor g218 (n_251, B[7], B[6]);
  nor g222 (n_290, B[5], B[6]);
  nand g223 (n_288, B[5], B[6]);
  xor g224 (n_252, B[7], A[0]);
  and g228 (n_423, A[0], n_249);
  xor g229 (n_257, B[7], A[1]);
  nand g230 (n_258, n_257, n_249);
  nand g231 (n_259, n_252, n_253);
  nand g232 (n_432, n_258, n_259);
  xor g233 (n_260, B[7], A[2]);
  nand g234 (n_261, n_260, n_249);
  nand g235 (n_262, n_257, n_253);
  nand g236 (n_439, n_261, n_262);
  xor g237 (n_263, B[7], A[3]);
  nand g238 (n_264, n_263, n_249);
  nand g239 (n_265, n_260, n_253);
  nand g240 (n_448, n_264, n_265);
  xor g241 (n_266, B[7], A[4]);
  nand g242 (n_267, n_266, n_249);
  nand g243 (n_268, n_263, n_253);
  nand g244 (n_457, n_267, n_268);
  xor g245 (n_269, B[7], A[5]);
  nand g246 (n_270, n_269, n_249);
  nand g247 (n_271, n_266, n_253);
  nand g248 (n_469, n_270, n_271);
  xor g249 (n_272, B[7], A[6]);
  nand g250 (n_273, n_272, n_249);
  nand g251 (n_274, n_269, n_253);
  nand g252 (n_483, n_273, n_274);
  xor g253 (n_275, B[7], A[7]);
  nand g254 (n_276, n_275, n_249);
  nand g255 (n_277, n_272, n_253);
  nand g256 (n_497, n_276, n_277);
  xor g257 (n_278, B[7], A[8]);
  nand g258 (n_279, n_278, n_249);
  nand g259 (n_280, n_275, n_253);
  nand g260 (n_514, n_279, n_280);
  xor g261 (n_281, B[7], A[9]);
  nand g262 (n_282, n_281, n_249);
  nand g263 (n_283, n_278, n_253);
  nand g264 (n_532, n_282, n_283);
  xor g265 (n_284, B[7], A[10]);
  nand g266 (n_285, n_284, n_249);
  nand g267 (n_286, n_281, n_253);
  nand g268 (n_552, n_285, n_286);
  or g271 (n_291, n_875, n_290);
  and g272 (n_428, B[7], n_291);
  xor g273 (n_292, B[8], B[7]);
  xor g274 (n_294, B[9], B[8]);
  nor g278 (n_327, B[7], B[8]);
  nand g279 (n_325, B[7], B[8]);
  xor g280 (n_295, B[9], A[0]);
  and g284 (n_437, A[0], n_292);
  xor g285 (n_300, B[9], A[1]);
  nand g286 (n_301, n_300, n_292);
  nand g287 (n_302, n_295, n_296);
  nand g288 (n_451, n_301, n_302);
  xor g289 (n_303, B[9], A[2]);
  nand g290 (n_304, n_303, n_292);
  nand g291 (n_305, n_300, n_296);
  nand g292 (n_462, n_304, n_305);
  xor g293 (n_306, B[9], A[3]);
  nand g294 (n_307, n_306, n_292);
  nand g295 (n_308, n_303, n_296);
  nand g296 (n_473, n_307, n_308);
  xor g297 (n_309, B[9], A[4]);
  nand g298 (n_310, n_309, n_292);
  nand g299 (n_311, n_306, n_296);
  nand g300 (n_488, n_310, n_311);
  xor g301 (n_312, B[9], A[5]);
  nand g302 (n_313, n_312, n_292);
  nand g303 (n_314, n_309, n_296);
  nand g304 (n_500, n_313, n_314);
  xor g305 (n_315, B[9], A[6]);
  nand g306 (n_316, n_315, n_292);
  nand g307 (n_317, n_312, n_296);
  nand g308 (n_517, n_316, n_317);
  xor g309 (n_318, B[9], A[7]);
  nand g310 (n_319, n_318, n_292);
  nand g311 (n_320, n_315, n_296);
  nand g312 (n_535, n_319, n_320);
  xor g313 (n_321, B[9], A[8]);
  nand g314 (n_322, n_321, n_292);
  nand g315 (n_323, n_318, n_296);
  nand g316 (n_555, n_322, n_323);
  or g319 (n_328, n_876, n_327);
  and g320 (n_447, B[9], n_328);
  xor g321 (n_329, B[10], B[9]);
  xor g322 (n_331, B[11], B[10]);
  nor g326 (n_358, B[9], B[10]);
  nand g327 (n_356, B[9], B[10]);
  xor g328 (n_332, B[11], A[0]);
  and g332 (n_459, A[0], n_329);
  xor g333 (n_337, B[11], A[1]);
  nand g334 (n_338, n_337, n_329);
  nand g335 (n_339, n_332, n_333);
  nand g336 (n_476, n_338, n_339);
  xor g337 (n_340, B[11], A[2]);
  nand g338 (n_341, n_340, n_329);
  nand g339 (n_342, n_337, n_333);
  nand g340 (n_489, n_341, n_342);
  xor g341 (n_343, B[11], A[3]);
  nand g342 (n_344, n_343, n_329);
  nand g343 (n_345, n_340, n_333);
  nand g344 (n_504, n_344, n_345);
  xor g345 (n_346, B[11], A[4]);
  nand g346 (n_347, n_346, n_329);
  nand g347 (n_348, n_343, n_333);
  nand g348 (n_521, n_347, n_348);
  xor g349 (n_349, B[11], A[5]);
  nand g350 (n_350, n_349, n_329);
  nand g351 (n_351, n_346, n_333);
  nand g352 (n_538, n_350, n_351);
  xor g353 (n_352, B[11], A[6]);
  nand g354 (n_353, n_352, n_329);
  nand g355 (n_354, n_349, n_333);
  nand g356 (n_558, n_353, n_354);
  or g359 (n_359, n_877, n_358);
  and g360 (n_470, B[11], n_359);
  xor g361 (n_360, B[12], B[11]);
  xor g362 (n_362, B[13], B[12]);
  nor g366 (n_383, B[11], B[12]);
  nand g367 (n_381, B[11], B[12]);
  xor g368 (n_363, B[13], A[0]);
  and g372 (n_485, A[0], n_360);
  xor g373 (n_368, B[13], A[1]);
  nand g374 (n_369, n_368, n_360);
  nand g375 (n_370, n_363, n_364);
  nand g376 (n_506, n_369, n_370);
  xor g377 (n_371, B[13], A[2]);
  nand g378 (n_372, n_371, n_360);
  nand g379 (n_373, n_368, n_364);
  nand g380 (n_522, n_372, n_373);
  xor g381 (n_374, B[13], A[3]);
  nand g382 (n_375, n_374, n_360);
  nand g383 (n_376, n_371, n_364);
  nand g384 (n_541, n_375, n_376);
  xor g385 (n_377, B[13], A[4]);
  nand g386 (n_378, n_377, n_360);
  nand g387 (n_379, n_374, n_364);
  nand g388 (n_561, n_378, n_379);
  or g391 (n_384, n_878, n_383);
  and g392 (n_499, B[13], n_384);
  xor g393 (n_385, B[14], B[13]);
  xor g394 (n_387, B[15], B[14]);
  nor g398 (n_402, B[13], B[14]);
  nand g399 (n_400, B[13], B[14]);
  xor g400 (n_388, B[15], A[0]);
  and g404 (n_516, A[0], n_385);
  xor g405 (n_393, B[15], A[1]);
  nand g406 (n_394, n_393, n_385);
  nand g407 (n_395, n_388, n_389);
  nand g408 (n_540, n_394, n_395);
  xor g409 (n_396, B[15], A[2]);
  nand g410 (n_397, n_396, n_385);
  nand g411 (n_398, n_393, n_389);
  nand g412 (n_559, n_397, n_398);
  or g415 (n_403, n_879, n_402);
  and g416 (n_534, B[15], n_403);
  and g428 (n_554, A[0], B[15]);
  xor g485 (n_80, n_412, n_413);
  and g486 (n_62, n_412, n_413);
  xor g487 (n_573, n_414, n_415);
  xor g488 (n_79, n_573, n_416);
  nand g489 (n_574, n_414, n_415);
  nand g490 (n_575, n_416, n_415);
  nand g491 (n_576, n_414, n_416);
  nand g492 (n_61, n_574, n_575, n_576);
  xor g493 (n_420, n_417, n_418);
  and g494 (n_424, n_417, n_418);
  xor g495 (n_577, n_419, n_420);
  xor g496 (n_78, n_577, n_421);
  nand g497 (n_578, n_419, n_420);
  nand g498 (n_579, n_421, n_420);
  nand g499 (n_580, n_419, n_421);
  nand g500 (n_60, n_578, n_579, n_580);
  xor g501 (n_581, n_422, n_423);
  xor g502 (n_427, n_581, n_424);
  nand g503 (n_582, n_422, n_423);
  nand g504 (n_583, n_424, n_423);
  nand g505 (n_584, n_422, n_424);
  nand g506 (n_434, n_582, n_583, n_584);
  xor g507 (n_585, n_425, n_426);
  xor g508 (n_77, n_585, n_427);
  nand g509 (n_586, n_425, n_426);
  nand g510 (n_587, n_427, n_426);
  nand g511 (n_588, n_425, n_427);
  nand g512 (n_59, n_586, n_587, n_588);
  xor g513 (n_433, n_428, n_429);
  and g514 (n_441, n_428, n_429);
  xor g515 (n_589, n_430, n_431);
  xor g516 (n_435, n_589, n_432);
  nand g517 (n_590, n_430, n_431);
  nand g518 (n_591, n_432, n_431);
  nand g519 (n_592, n_430, n_432);
  nand g520 (n_443, n_590, n_591, n_592);
  xor g521 (n_593, n_433, n_434);
  xor g522 (n_76, n_593, n_435);
  nand g523 (n_594, n_433, n_434);
  nand g524 (n_595, n_435, n_434);
  nand g525 (n_596, n_433, n_435);
  nand g526 (n_58, n_594, n_595, n_596);
  xor g527 (n_597, n_436, n_437);
  xor g528 (n_442, n_597, n_438);
  nand g529 (n_598, n_436, n_437);
  nand g530 (n_599, n_438, n_437);
  nand g531 (n_600, n_436, n_438);
  nand g532 (n_452, n_598, n_599, n_600);
  xor g533 (n_601, n_439, n_440);
  xor g534 (n_444, n_601, n_441);
  nand g535 (n_602, n_439, n_440);
  nand g536 (n_603, n_441, n_440);
  nand g537 (n_604, n_439, n_441);
  nand g538 (n_453, n_602, n_603, n_604);
  xor g539 (n_605, n_442, n_443);
  xor g540 (n_75, n_605, n_444);
  nand g541 (n_606, n_442, n_443);
  nand g542 (n_607, n_444, n_443);
  nand g543 (n_608, n_442, n_444);
  nand g544 (n_57, n_606, n_607, n_608);
  xor g545 (n_449, n_445, n_446);
  and g546 (n_461, n_445, n_446);
  xor g547 (n_609, n_447, n_448);
  xor g548 (n_454, n_609, n_449);
  nand g549 (n_610, n_447, n_448);
  nand g550 (n_611, n_449, n_448);
  nand g551 (n_612, n_447, n_449);
  nand g552 (n_463, n_610, n_611, n_612);
  xor g553 (n_613, n_450, n_451);
  xor g554 (n_455, n_613, n_452);
  nand g555 (n_614, n_450, n_451);
  nand g556 (n_615, n_452, n_451);
  nand g557 (n_616, n_450, n_452);
  nand g558 (n_466, n_614, n_615, n_616);
  xor g559 (n_617, n_453, n_454);
  xor g560 (n_74, n_617, n_455);
  nand g561 (n_618, n_453, n_454);
  nand g562 (n_619, n_455, n_454);
  nand g563 (n_620, n_453, n_455);
  nand g564 (n_56, n_618, n_619, n_620);
  xor g565 (n_621, n_456, n_457);
  xor g566 (n_464, n_621, n_458);
  nand g567 (n_622, n_456, n_457);
  nand g568 (n_623, n_458, n_457);
  nand g569 (n_624, n_456, n_458);
  nand g570 (n_475, n_622, n_623, n_624);
  xor g571 (n_625, n_459, n_460);
  xor g572 (n_465, n_625, n_461);
  nand g573 (n_626, n_459, n_460);
  nand g574 (n_627, n_461, n_460);
  nand g575 (n_628, n_459, n_461);
  nand g576 (n_477, n_626, n_627, n_628);
  xor g577 (n_629, n_462, n_463);
  xor g578 (n_467, n_629, n_464);
  nand g579 (n_630, n_462, n_463);
  nand g580 (n_631, n_464, n_463);
  nand g581 (n_632, n_462, n_464);
  nand g582 (n_480, n_630, n_631, n_632);
  xor g583 (n_633, n_465, n_466);
  xor g584 (n_73, n_633, n_467);
  nand g585 (n_634, n_465, n_466);
  nand g586 (n_635, n_467, n_466);
  nand g587 (n_636, n_465, n_467);
  nand g588 (n_55, n_634, n_635, n_636);
  xor g589 (n_474, n_468, n_469);
  and g590 (n_487, n_468, n_469);
  xor g591 (n_637, n_470, n_471);
  xor g592 (n_478, n_637, n_472);
  nand g593 (n_638, n_470, n_471);
  nand g594 (n_639, n_472, n_471);
  nand g595 (n_640, n_470, n_472);
  nand g596 (n_491, n_638, n_639, n_640);
  xor g597 (n_641, n_473, n_474);
  xor g598 (n_479, n_641, n_475);
  nand g599 (n_642, n_473, n_474);
  nand g600 (n_643, n_475, n_474);
  nand g601 (n_644, n_473, n_475);
  nand g602 (n_493, n_642, n_643, n_644);
  xor g603 (n_645, n_476, n_477);
  xor g604 (n_481, n_645, n_478);
  nand g605 (n_646, n_476, n_477);
  nand g606 (n_647, n_478, n_477);
  nand g607 (n_648, n_476, n_478);
  nand g608 (n_495, n_646, n_647, n_648);
  xor g609 (n_649, n_479, n_480);
  xor g610 (n_72, n_649, n_481);
  nand g611 (n_650, n_479, n_480);
  nand g612 (n_651, n_481, n_480);
  nand g613 (n_652, n_479, n_481);
  nand g614 (n_54, n_650, n_651, n_652);
  xor g615 (n_653, n_482, n_483);
  xor g616 (n_490, n_653, n_484);
  nand g617 (n_654, n_482, n_483);
  nand g618 (n_655, n_484, n_483);
  nand g619 (n_656, n_482, n_484);
  nand g620 (n_505, n_654, n_655, n_656);
  xor g621 (n_657, n_485, n_486);
  xor g622 (n_492, n_657, n_487);
  nand g623 (n_658, n_485, n_486);
  nand g624 (n_659, n_487, n_486);
  nand g625 (n_660, n_485, n_487);
  nand g626 (n_507, n_658, n_659, n_660);
  xor g627 (n_661, n_488, n_489);
  xor g628 (n_494, n_661, n_490);
  nand g629 (n_662, n_488, n_489);
  nand g630 (n_663, n_490, n_489);
  nand g631 (n_664, n_488, n_490);
  nand g632 (n_509, n_662, n_663, n_664);
  xor g633 (n_665, n_491, n_492);
  xor g634 (n_496, n_665, n_493);
  nand g635 (n_666, n_491, n_492);
  nand g636 (n_667, n_493, n_492);
  nand g637 (n_668, n_491, n_493);
  nand g638 (n_512, n_666, n_667, n_668);
  xor g639 (n_669, n_494, n_495);
  xor g640 (n_71, n_669, n_496);
  nand g641 (n_670, n_494, n_495);
  nand g642 (n_671, n_496, n_495);
  nand g643 (n_672, n_494, n_496);
  nand g644 (n_53, n_670, n_671, n_672);
  xor g645 (n_502, n_497, n_498);
  and g646 (n_520, n_497, n_498);
  xor g647 (n_673, n_499, n_500);
  xor g648 (n_508, n_673, n_501);
  nand g649 (n_674, n_499, n_500);
  nand g650 (n_675, n_501, n_500);
  nand g651 (n_676, n_499, n_501);
  nand g652 (n_523, n_674, n_675, n_676);
  xor g653 (n_677, n_502, n_503);
  xor g654 (n_510, n_677, n_504);
  nand g655 (n_678, n_502, n_503);
  nand g656 (n_679, n_504, n_503);
  nand g657 (n_680, n_502, n_504);
  nand g658 (n_525, n_678, n_679, n_680);
  xor g659 (n_681, n_505, n_506);
  xor g660 (n_511, n_681, n_507);
  nand g661 (n_682, n_505, n_506);
  nand g662 (n_683, n_507, n_506);
  nand g663 (n_684, n_505, n_507);
  nand g664 (n_528, n_682, n_683, n_684);
  xor g665 (n_685, n_508, n_509);
  xor g666 (n_513, n_685, n_510);
  nand g667 (n_686, n_508, n_509);
  nand g668 (n_687, n_510, n_509);
  nand g669 (n_688, n_508, n_510);
  nand g670 (n_530, n_686, n_687, n_688);
  xor g671 (n_689, n_511, n_512);
  xor g672 (n_70, n_689, n_513);
  nand g673 (n_690, n_511, n_512);
  nand g674 (n_691, n_513, n_512);
  nand g675 (n_692, n_511, n_513);
  nand g676 (n_52, n_690, n_691, n_692);
  xor g677 (n_693, n_514, n_515);
  xor g678 (n_524, n_693, n_516);
  nand g679 (n_694, n_514, n_515);
  nand g680 (n_695, n_516, n_515);
  nand g681 (n_696, n_514, n_516);
  nand g682 (n_542, n_694, n_695, n_696);
  xor g683 (n_697, n_517, n_518);
  xor g684 (n_526, n_697, n_519);
  nand g685 (n_698, n_517, n_518);
  nand g686 (n_699, n_519, n_518);
  nand g687 (n_700, n_517, n_519);
  nand g688 (n_543, n_698, n_699, n_700);
  xor g689 (n_701, n_520, n_521);
  xor g690 (n_527, n_701, n_522);
  nand g691 (n_702, n_520, n_521);
  nand g692 (n_703, n_522, n_521);
  nand g693 (n_704, n_520, n_522);
  nand g694 (n_546, n_702, n_703, n_704);
  xor g695 (n_705, n_523, n_524);
  xor g696 (n_529, n_705, n_525);
  nand g697 (n_706, n_523, n_524);
  nand g698 (n_707, n_525, n_524);
  nand g699 (n_708, n_523, n_525);
  nand g700 (n_548, n_706, n_707, n_708);
  xor g701 (n_709, n_526, n_527);
  xor g702 (n_531, n_709, n_528);
  nand g703 (n_710, n_526, n_527);
  nand g704 (n_711, n_528, n_527);
  nand g705 (n_712, n_526, n_528);
  nand g706 (n_550, n_710, n_711, n_712);
  xor g707 (n_713, n_529, n_530);
  xor g708 (n_69, n_713, n_531);
  nand g709 (n_714, n_529, n_530);
  nand g710 (n_715, n_531, n_530);
  nand g711 (n_716, n_529, n_531);
  nand g712 (n_51, n_714, n_715, n_716);
  xor g713 (n_539, n_532, n_533);
  and g714 (n_560, n_532, n_533);
  xor g715 (n_717, n_534, n_535);
  xor g716 (n_544, n_717, n_536);
  nand g717 (n_718, n_534, n_535);
  nand g718 (n_719, n_536, n_535);
  nand g719 (n_720, n_534, n_536);
  nand g720 (n_563, n_718, n_719, n_720);
  xor g721 (n_721, n_537, n_538);
  xor g722 (n_545, n_721, n_539);
  nand g723 (n_722, n_537, n_538);
  nand g724 (n_723, n_539, n_538);
  nand g725 (n_724, n_537, n_539);
  nand g726 (n_565, n_722, n_723, n_724);
  xor g727 (n_725, n_540, n_541);
  xor g728 (n_547, n_725, n_542);
  nand g729 (n_726, n_540, n_541);
  nand g730 (n_727, n_542, n_541);
  nand g731 (n_728, n_540, n_542);
  nand g732 (n_567, n_726, n_727, n_728);
  xor g733 (n_729, n_543, n_544);
  xor g734 (n_549, n_729, n_545);
  nand g735 (n_730, n_543, n_544);
  nand g736 (n_731, n_545, n_544);
  nand g737 (n_732, n_543, n_545);
  nand g738 (n_569, n_730, n_731, n_732);
  xor g739 (n_733, n_546, n_547);
  xor g740 (n_551, n_733, n_548);
  nand g741 (n_734, n_546, n_547);
  nand g742 (n_735, n_548, n_547);
  nand g743 (n_736, n_546, n_548);
  nand g744 (n_571, n_734, n_735, n_736);
  xor g745 (n_737, n_549, n_550);
  xor g746 (n_68, n_737, n_551);
  nand g747 (n_738, n_549, n_550);
  nand g748 (n_739, n_551, n_550);
  nand g749 (n_740, n_549, n_551);
  nand g750 (n_50, n_738, n_739, n_740);
  xor g751 (n_741, n_552, n_553);
  xor g752 (n_562, n_741, n_554);
  xor g757 (n_745, n_555, n_556);
  xor g758 (n_564, n_745, n_557);
  xor g763 (n_749, n_558, n_559);
  xor g764 (n_566, n_749, n_560);
  xor g769 (n_753, n_561, n_562);
  xor g770 (n_568, n_753, n_563);
  xor g775 (n_757, n_564, n_565);
  xor g776 (n_570, n_757, n_566);
  xor g781 (n_761, n_567, n_568);
  xor g782 (n_572, n_761, n_569);
  xor g787 (n_765, n_570, n_571);
  xor g788 (n_67, n_765, n_572);
  nor g800 (n_774, n_65, n_82);
  nand g801 (n_777, n_65, n_82);
  nor g802 (n_779, n_64, n_81);
  nand g803 (n_782, n_64, n_81);
  nor g804 (n_784, n_63, n_80);
  nand g805 (n_787, n_63, n_80);
  nor g806 (n_789, n_62, n_79);
  nand g807 (n_792, n_62, n_79);
  nor g808 (n_794, n_61, n_78);
  nand g809 (n_797, n_61, n_78);
  nor g810 (n_799, n_60, n_77);
  nand g811 (n_802, n_60, n_77);
  nor g812 (n_804, n_59, n_76);
  nand g813 (n_807, n_59, n_76);
  nor g814 (n_809, n_58, n_75);
  nand g815 (n_812, n_58, n_75);
  nor g816 (n_814, n_57, n_74);
  nand g817 (n_817, n_57, n_74);
  nor g818 (n_819, n_56, n_73);
  nand g819 (n_822, n_56, n_73);
  nor g820 (n_824, n_55, n_72);
  nand g821 (n_827, n_55, n_72);
  nor g822 (n_829, n_54, n_71);
  nand g823 (n_832, n_54, n_71);
  nor g824 (n_834, n_53, n_70);
  nand g825 (n_837, n_53, n_70);
  nor g826 (n_839, n_52, n_69);
  nand g827 (n_842, n_52, n_69);
  nor g828 (n_844, n_51, n_68);
  nand g829 (n_847, n_51, n_68);
  nand g837 (n_785, n_782, n_886);
  nand g840 (n_790, n_787, n_891);
  nand g843 (n_795, n_792, n_895);
  nand g846 (n_800, n_797, n_901);
  nand g849 (n_805, n_802, n_905);
  nand g852 (n_810, n_807, n_907);
  nand g855 (n_815, n_812, n_908);
  nand g858 (n_820, n_817, n_909);
  nand g861 (n_825, n_822, n_910);
  nand g864 (n_830, n_827, n_911);
  nand g867 (n_835, n_832, n_912);
  nand g870 (n_840, n_837, n_913);
  nand g873 (n_845, n_842, n_914);
  nand g876 (n_850, n_847, n_915);
  xnor g883 (Z[3], n_785, n_885);
  xnor g885 (Z[4], n_790, n_888);
  xnor g887 (Z[5], n_795, n_889);
  xnor g889 (Z[6], n_800, n_890);
  xnor g891 (Z[7], n_805, n_892);
  xnor g893 (Z[8], n_810, n_893);
  xnor g895 (Z[9], n_815, n_894);
  xnor g897 (Z[10], n_820, n_896);
  xnor g899 (Z[11], n_825, n_897);
  xnor g901 (Z[12], n_830, n_898);
  xnor g903 (Z[13], n_835, n_902);
  xnor g905 (Z[14], n_840, n_903);
  xnor g907 (Z[15], n_845, n_904);
  xnor g909 (Z[16], n_850, n_906);
  and g912 (n_873, wc, n_196);
  not gc (wc, A[0]);
  and g913 (n_874, wc0, n_245);
  not gc0 (wc0, A[0]);
  and g914 (n_875, wc1, n_288);
  not gc1 (wc1, A[0]);
  and g915 (n_876, wc2, n_325);
  not gc2 (wc2, A[0]);
  and g916 (n_877, wc3, n_356);
  not gc3 (wc3, A[0]);
  and g917 (n_878, wc4, n_381);
  not gc4 (wc4, A[0]);
  and g918 (n_879, wc5, n_400);
  not gc5 (wc5, A[0]);
  and g919 (n_89, wc6, n_87);
  not gc6 (wc6, B[0]);
  and g921 (n_149, n_147, wc7);
  not gc7 (wc7, n_145);
  and g922 (n_204, n_202, wc8);
  not gc8 (wc8, n_200);
  and g923 (n_253, n_251, wc9);
  not gc9 (wc9, n_249);
  and g924 (n_296, n_294, wc10);
  not gc10 (wc10, n_292);
  and g925 (n_333, n_331, wc11);
  not gc11 (wc11, n_329);
  and g926 (n_364, n_362, wc12);
  not gc12 (wc12, n_360);
  and g927 (n_389, n_387, wc13);
  not gc13 (wc13, n_385);
  and g928 (n_65, B[1], wc14);
  not gc14 (wc14, Z[0]);
  or g929 (n_882, wc15, n_774);
  not gc15 (wc15, n_777);
  or g930 (n_883, wc16, n_779);
  not gc16 (wc16, n_782);
  not g932 (Z[1], n_882);
  or g933 (n_885, wc17, n_784);
  not gc17 (wc17, n_787);
  or g934 (n_886, n_777, n_779);
  xor g935 (Z[2], n_777, n_883);
  or g936 (n_888, wc18, n_789);
  not gc18 (wc18, n_792);
  or g937 (n_889, wc19, n_794);
  not gc19 (wc19, n_797);
  or g938 (n_890, wc20, n_799);
  not gc20 (wc20, n_802);
  or g939 (n_891, wc21, n_784);
  not gc21 (wc21, n_785);
  or g940 (n_892, wc22, n_804);
  not gc22 (wc22, n_807);
  or g941 (n_893, wc23, n_809);
  not gc23 (wc23, n_812);
  or g942 (n_894, wc24, n_814);
  not gc24 (wc24, n_817);
  or g943 (n_895, wc25, n_789);
  not gc25 (wc25, n_790);
  or g944 (n_896, wc26, n_819);
  not gc26 (wc26, n_822);
  or g945 (n_897, wc27, n_824);
  not gc27 (wc27, n_827);
  or g946 (n_898, wc28, n_829);
  not gc28 (wc28, n_832);
  and g947 (n_899, n_50, n_67);
  or g948 (n_900, n_50, n_67);
  or g949 (n_901, wc29, n_794);
  not gc29 (wc29, n_795);
  or g950 (n_902, wc30, n_834);
  not gc30 (wc30, n_837);
  or g951 (n_903, wc31, n_839);
  not gc31 (wc31, n_842);
  or g952 (n_904, wc32, n_844);
  not gc32 (wc32, n_847);
  or g953 (n_905, wc33, n_799);
  not gc33 (wc33, n_800);
  or g954 (n_906, wc34, n_899);
  not gc34 (wc34, n_900);
  or g955 (n_907, wc35, n_804);
  not gc35 (wc35, n_805);
  or g956 (n_908, wc36, n_809);
  not gc36 (wc36, n_810);
  or g957 (n_909, wc37, n_814);
  not gc37 (wc37, n_815);
  or g958 (n_910, wc38, n_819);
  not gc38 (wc38, n_820);
  or g959 (n_911, wc39, n_824);
  not gc39 (wc39, n_825);
  or g960 (n_912, wc40, n_829);
  not gc40 (wc40, n_830);
  or g961 (n_913, wc41, n_834);
  not gc41 (wc41, n_835);
  or g962 (n_914, wc42, n_839);
  not gc42 (wc42, n_840);
  or g963 (n_915, wc43, n_844);
  not gc43 (wc43, n_845);
endmodule

module mult_unsigned_120_GENERIC(A, B, Z);
  input [15:0] A, B;
  output [16:0] Z;
  wire [15:0] A, B;
  wire [16:0] Z;
  mult_unsigned_120_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module mult_unsigned_35_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $unsigned(A) * $unsigned(B);"
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_325;
  wire n_328, n_330, n_333, n_335, n_336, n_338, n_340, n_341;
  wire n_343, n_345, n_346, n_348, n_350, n_351, n_353, n_355;
  wire n_356, n_358, n_360, n_361, n_363, n_365, n_366, n_368;
  wire n_370, n_371, n_373, n_375, n_376, n_378, n_380, n_381;
  wire n_383, n_385, n_386, n_388, n_390, n_391, n_393, n_417;
  wire n_419, n_420, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445;
  and g1 (Z[0], A[0], B[0]);
  and g2 (n_46, A[1], B[0]);
  and g3 (n_63, A[2], B[0]);
  and g4 (n_67, A[3], B[0]);
  and g5 (n_72, A[4], B[0]);
  and g6 (n_80, A[5], B[0]);
  and g7 (n_90, A[6], B[0]);
  and g8 (n_103, A[7], B[0]);
  and g9 (n_61, A[0], B[1]);
  and g10 (n_45, A[1], B[1]);
  and g11 (n_68, A[2], B[1]);
  and g12 (n_73, A[3], B[1]);
  and g13 (n_64, A[4], B[1]);
  and g14 (n_91, A[5], B[1]);
  and g15 (n_104, A[6], B[1]);
  and g16 (n_120, A[7], B[1]);
  and g17 (n_66, A[0], B[2]);
  and g18 (n_70, A[1], B[2]);
  and g19 (n_76, A[2], B[2]);
  and g20 (n_83, A[3], B[2]);
  and g21 (n_94, A[4], B[2]);
  and g22 (n_108, A[5], B[2]);
  and g23 (n_121, A[6], B[2]);
  and g24 (n_137, A[7], B[2]);
  and g25 (n_69, A[0], B[3]);
  and g26 (n_74, A[1], B[3]);
  and g27 (n_81, A[2], B[3]);
  and g28 (n_92, A[3], B[3]);
  and g29 (n_105, A[4], B[3]);
  and g30 (n_124, A[5], B[3]);
  and g31 (n_138, A[6], B[3]);
  and g32 (n_152, A[7], B[3]);
  and g33 (n_75, A[0], B[4]);
  and g34 (n_82, A[1], B[4]);
  and g35 (n_93, A[2], B[4]);
  and g36 (n_107, A[3], B[4]);
  and g37 (n_122, A[4], B[4]);
  and g38 (n_141, A[5], B[4]);
  and g39 (n_153, A[6], B[4]);
  and g40 (n_164, A[7], B[4]);
  and g41 (n_84, A[0], B[5]);
  and g42 (n_65, A[1], B[5]);
  and g43 (n_109, A[2], B[5]);
  and g44 (n_123, A[3], B[5]);
  and g45 (n_139, A[4], B[5]);
  and g46 (n_156, A[5], B[5]);
  and g47 (n_165, A[6], B[5]);
  and g48 (n_173, A[7], B[5]);
  and g49 (n_95, A[0], B[6]);
  and g50 (n_110, A[1], B[6]);
  and g51 (n_125, A[2], B[6]);
  and g52 (n_140, A[3], B[6]);
  and g53 (n_154, A[4], B[6]);
  and g54 (n_167, A[5], B[6]);
  and g55 (n_174, A[6], B[6]);
  and g56 (n_179, A[7], B[6]);
  and g57 (n_106, A[0], B[7]);
  and g58 (n_126, A[1], B[7]);
  and g59 (n_142, A[2], B[7]);
  and g60 (n_155, A[3], B[7]);
  and g61 (n_166, A[4], B[7]);
  and g62 (n_175, A[5], B[7]);
  and g63 (n_180, A[6], B[7]);
  and g64 (n_33, A[7], B[7]);
  xor g107 (n_60, n_63, n_66);
  and g108 (n_44, n_63, n_66);
  xor g109 (n_71, n_67, n_68);
  and g110 (n_78, n_67, n_68);
  xor g111 (n_182, n_69, n_70);
  xor g112 (n_59, n_182, n_71);
  nand g113 (n_183, n_69, n_70);
  nand g114 (n_184, n_71, n_70);
  nand g115 (n_185, n_69, n_71);
  nand g116 (n_43, n_183, n_184, n_185);
  xor g117 (n_77, n_72, n_73);
  and g118 (n_86, n_72, n_73);
  xor g119 (n_186, n_74, n_75);
  xor g120 (n_79, n_186, n_76);
  nand g121 (n_187, n_74, n_75);
  nand g122 (n_188, n_76, n_75);
  nand g123 (n_189, n_74, n_76);
  nand g124 (n_87, n_187, n_188, n_189);
  xor g125 (n_190, n_77, n_78);
  xor g126 (n_58, n_190, n_79);
  nand g127 (n_191, n_77, n_78);
  nand g128 (n_192, n_79, n_78);
  nand g129 (n_193, n_77, n_79);
  nand g130 (n_42, n_191, n_192, n_193);
  xor g131 (n_85, n_80, n_64);
  and g132 (n_96, n_80, n_64);
  xor g133 (n_194, n_81, n_82);
  xor g134 (n_88, n_194, n_83);
  nand g135 (n_195, n_81, n_82);
  nand g136 (n_196, n_83, n_82);
  nand g137 (n_197, n_81, n_83);
  nand g138 (n_98, n_195, n_196, n_197);
  xor g139 (n_198, n_84, n_85);
  xor g140 (n_89, n_198, n_86);
  nand g141 (n_199, n_84, n_85);
  nand g142 (n_200, n_86, n_85);
  nand g143 (n_201, n_84, n_86);
  nand g144 (n_100, n_199, n_200, n_201);
  xor g145 (n_202, n_87, n_88);
  xor g146 (n_57, n_202, n_89);
  nand g147 (n_203, n_87, n_88);
  nand g148 (n_204, n_89, n_88);
  nand g149 (n_205, n_87, n_89);
  nand g150 (n_41, n_203, n_204, n_205);
  xor g151 (n_97, n_90, n_91);
  and g152 (n_111, n_90, n_91);
  xor g153 (n_206, n_92, n_93);
  xor g154 (n_99, n_206, n_94);
  nand g155 (n_207, n_92, n_93);
  nand g156 (n_208, n_94, n_93);
  nand g157 (n_209, n_92, n_94);
  nand g158 (n_113, n_207, n_208, n_209);
  xor g159 (n_210, n_65, n_95);
  xor g160 (n_101, n_210, n_96);
  nand g161 (n_211, n_65, n_95);
  nand g162 (n_212, n_96, n_95);
  nand g163 (n_213, n_65, n_96);
  nand g164 (n_116, n_211, n_212, n_213);
  xor g165 (n_214, n_97, n_98);
  xor g166 (n_102, n_214, n_99);
  nand g167 (n_215, n_97, n_98);
  nand g168 (n_216, n_99, n_98);
  nand g169 (n_217, n_97, n_99);
  nand g170 (n_118, n_215, n_216, n_217);
  xor g171 (n_218, n_100, n_101);
  xor g172 (n_56, n_218, n_102);
  nand g173 (n_219, n_100, n_101);
  nand g174 (n_220, n_102, n_101);
  nand g175 (n_221, n_100, n_102);
  nand g176 (n_40, n_219, n_220, n_221);
  xor g177 (n_112, n_103, n_104);
  and g178 (n_128, n_103, n_104);
  xor g179 (n_222, n_105, n_106);
  xor g180 (n_115, n_222, n_107);
  nand g181 (n_223, n_105, n_106);
  nand g182 (n_224, n_107, n_106);
  nand g183 (n_225, n_105, n_107);
  nand g184 (n_129, n_223, n_224, n_225);
  xor g185 (n_226, n_108, n_109);
  xor g186 (n_114, n_226, n_110);
  nand g187 (n_227, n_108, n_109);
  nand g188 (n_228, n_110, n_109);
  nand g189 (n_229, n_108, n_110);
  nand g190 (n_130, n_227, n_228, n_229);
  xor g191 (n_230, n_111, n_112);
  xor g192 (n_117, n_230, n_113);
  nand g193 (n_231, n_111, n_112);
  nand g194 (n_232, n_113, n_112);
  nand g195 (n_233, n_111, n_113);
  nand g196 (n_133, n_231, n_232, n_233);
  xor g197 (n_234, n_114, n_115);
  xor g198 (n_119, n_234, n_116);
  nand g199 (n_235, n_114, n_115);
  nand g200 (n_236, n_116, n_115);
  nand g201 (n_237, n_114, n_116);
  nand g202 (n_135, n_235, n_236, n_237);
  xor g203 (n_238, n_117, n_118);
  xor g204 (n_55, n_238, n_119);
  nand g205 (n_239, n_117, n_118);
  nand g206 (n_240, n_119, n_118);
  nand g207 (n_241, n_117, n_119);
  nand g208 (n_39, n_239, n_240, n_241);
  xor g209 (n_127, n_120, n_121);
  and g210 (n_143, n_120, n_121);
  xor g211 (n_242, n_122, n_123);
  xor g212 (n_131, n_242, n_124);
  nand g213 (n_243, n_122, n_123);
  nand g214 (n_244, n_124, n_123);
  nand g215 (n_245, n_122, n_124);
  nand g216 (n_144, n_243, n_244, n_245);
  xor g217 (n_246, n_125, n_126);
  xor g218 (n_132, n_246, n_127);
  nand g219 (n_247, n_125, n_126);
  nand g220 (n_248, n_127, n_126);
  nand g221 (n_249, n_125, n_127);
  nand g222 (n_147, n_247, n_248, n_249);
  xor g223 (n_250, n_128, n_129);
  xor g224 (n_134, n_250, n_130);
  nand g225 (n_251, n_128, n_129);
  nand g226 (n_252, n_130, n_129);
  nand g227 (n_253, n_128, n_130);
  nand g228 (n_148, n_251, n_252, n_253);
  xor g229 (n_254, n_131, n_132);
  xor g230 (n_136, n_254, n_133);
  nand g231 (n_255, n_131, n_132);
  nand g232 (n_256, n_133, n_132);
  nand g233 (n_257, n_131, n_133);
  nand g234 (n_151, n_255, n_256, n_257);
  xor g235 (n_258, n_134, n_135);
  xor g236 (n_54, n_258, n_136);
  nand g237 (n_259, n_134, n_135);
  nand g238 (n_260, n_136, n_135);
  nand g239 (n_261, n_134, n_136);
  nand g240 (n_38, n_259, n_260, n_261);
  xor g241 (n_262, n_137, n_138);
  xor g242 (n_146, n_262, n_139);
  nand g243 (n_263, n_137, n_138);
  nand g244 (n_264, n_139, n_138);
  nand g245 (n_265, n_137, n_139);
  nand g246 (n_158, n_263, n_264, n_265);
  xor g247 (n_266, n_140, n_141);
  xor g248 (n_145, n_266, n_142);
  nand g249 (n_267, n_140, n_141);
  nand g250 (n_268, n_142, n_141);
  nand g251 (n_269, n_140, n_142);
  nand g252 (n_157, n_267, n_268, n_269);
  xor g253 (n_270, n_143, n_144);
  xor g254 (n_149, n_270, n_145);
  nand g255 (n_271, n_143, n_144);
  nand g256 (n_272, n_145, n_144);
  nand g257 (n_273, n_143, n_145);
  nand g258 (n_161, n_271, n_272, n_273);
  xor g259 (n_274, n_146, n_147);
  xor g260 (n_150, n_274, n_148);
  nand g261 (n_275, n_146, n_147);
  nand g262 (n_276, n_148, n_147);
  nand g263 (n_277, n_146, n_148);
  nand g264 (n_163, n_275, n_276, n_277);
  xor g265 (n_278, n_149, n_150);
  xor g266 (n_53, n_278, n_151);
  nand g267 (n_279, n_149, n_150);
  nand g268 (n_280, n_151, n_150);
  nand g269 (n_281, n_149, n_151);
  nand g270 (n_37, n_279, n_280, n_281);
  xor g271 (n_282, n_152, n_153);
  xor g272 (n_159, n_282, n_154);
  nand g273 (n_283, n_152, n_153);
  nand g274 (n_284, n_154, n_153);
  nand g275 (n_285, n_152, n_154);
  nand g276 (n_168, n_283, n_284, n_285);
  xor g277 (n_286, n_155, n_156);
  xor g278 (n_160, n_286, n_157);
  nand g279 (n_287, n_155, n_156);
  nand g280 (n_288, n_157, n_156);
  nand g281 (n_289, n_155, n_157);
  nand g282 (n_170, n_287, n_288, n_289);
  xor g283 (n_290, n_158, n_159);
  xor g284 (n_162, n_290, n_160);
  nand g285 (n_291, n_158, n_159);
  nand g286 (n_292, n_160, n_159);
  nand g287 (n_293, n_158, n_160);
  nand g288 (n_172, n_291, n_292, n_293);
  xor g289 (n_294, n_161, n_162);
  xor g290 (n_52, n_294, n_163);
  nand g291 (n_295, n_161, n_162);
  nand g292 (n_296, n_163, n_162);
  nand g293 (n_297, n_161, n_163);
  nand g294 (n_36, n_295, n_296, n_297);
  xor g295 (n_298, n_164, n_165);
  xor g296 (n_169, n_298, n_166);
  nand g297 (n_299, n_164, n_165);
  nand g298 (n_300, n_166, n_165);
  nand g299 (n_301, n_164, n_166);
  nand g300 (n_176, n_299, n_300, n_301);
  xor g301 (n_302, n_167, n_168);
  xor g302 (n_171, n_302, n_169);
  nand g303 (n_303, n_167, n_168);
  nand g304 (n_304, n_169, n_168);
  nand g305 (n_305, n_167, n_169);
  nand g306 (n_178, n_303, n_304, n_305);
  xor g307 (n_306, n_170, n_171);
  xor g308 (n_51, n_306, n_172);
  nand g309 (n_307, n_170, n_171);
  nand g310 (n_308, n_172, n_171);
  nand g311 (n_309, n_170, n_172);
  nand g312 (n_50, n_307, n_308, n_309);
  xor g313 (n_310, n_173, n_174);
  xor g314 (n_177, n_310, n_175);
  nand g315 (n_311, n_173, n_174);
  nand g316 (n_312, n_175, n_174);
  nand g317 (n_313, n_173, n_175);
  nand g318 (n_181, n_311, n_312, n_313);
  xor g319 (n_314, n_176, n_177);
  xor g320 (n_35, n_314, n_178);
  nand g321 (n_315, n_176, n_177);
  nand g322 (n_316, n_178, n_177);
  nand g323 (n_317, n_176, n_178);
  nand g324 (n_49, n_315, n_316, n_317);
  xor g325 (n_318, n_179, n_180);
  xor g326 (n_34, n_318, n_181);
  nand g327 (n_319, n_179, n_180);
  nand g328 (n_320, n_181, n_180);
  nand g329 (n_321, n_179, n_181);
  nand g330 (n_48, n_319, n_320, n_321);
  nor g336 (n_325, n_46, n_61);
  nand g337 (n_328, n_46, n_61);
  nor g338 (n_330, n_45, n_60);
  nand g339 (n_333, n_45, n_60);
  nor g340 (n_335, n_44, n_59);
  nand g341 (n_338, n_44, n_59);
  nor g342 (n_340, n_43, n_58);
  nand g343 (n_343, n_43, n_58);
  nor g344 (n_345, n_42, n_57);
  nand g345 (n_348, n_42, n_57);
  nor g346 (n_350, n_41, n_56);
  nand g347 (n_353, n_41, n_56);
  nor g348 (n_355, n_40, n_55);
  nand g349 (n_358, n_40, n_55);
  nor g350 (n_360, n_39, n_54);
  nand g351 (n_363, n_39, n_54);
  nor g352 (n_365, n_38, n_53);
  nand g353 (n_368, n_38, n_53);
  nor g354 (n_370, n_37, n_52);
  nand g355 (n_373, n_37, n_52);
  nor g356 (n_375, n_36, n_51);
  nand g357 (n_378, n_36, n_51);
  nor g358 (n_380, n_35, n_50);
  nand g359 (n_383, n_35, n_50);
  nor g360 (n_385, n_34, n_49);
  nand g361 (n_388, n_34, n_49);
  nor g362 (n_390, n_33, n_48);
  nand g363 (n_393, n_33, n_48);
  nand g371 (n_336, n_333, n_420);
  nand g374 (n_341, n_338, n_424);
  nand g377 (n_346, n_343, n_428);
  nand g380 (n_351, n_348, n_434);
  nand g383 (n_356, n_353, n_437);
  nand g386 (n_361, n_358, n_438);
  nand g389 (n_366, n_363, n_439);
  nand g392 (n_371, n_368, n_440);
  nand g65 (n_376, n_373, n_441);
  nand g68 (n_381, n_378, n_442);
  nand g71 (n_386, n_383, n_443);
  nand g74 (n_391, n_388, n_444);
  nand g77 (Z[15], n_393, n_445);
  xnor g86 (Z[3], n_336, n_422);
  xnor g88 (Z[4], n_341, n_423);
  xnor g90 (Z[5], n_346, n_425);
  xnor g92 (Z[6], n_351, n_427);
  xnor g94 (Z[7], n_356, n_429);
  xnor g96 (Z[8], n_361, n_431);
  xnor g98 (Z[9], n_366, n_432);
  xnor g100 (Z[10], n_371, n_435);
  xnor g102 (Z[11], n_376, n_436);
  xnor g104 (Z[12], n_381, n_433);
  xnor g106 (Z[13], n_386, n_430);
  xnor g396 (Z[14], n_391, n_426);
  or g400 (n_417, wc, n_325);
  not gc (wc, n_328);
  not g402 (Z[1], n_417);
  or g403 (n_419, wc0, n_330);
  not gc0 (wc0, n_333);
  or g404 (n_420, n_328, n_330);
  xor g405 (Z[2], n_328, n_419);
  or g406 (n_422, wc1, n_335);
  not gc1 (wc1, n_338);
  or g407 (n_423, wc2, n_340);
  not gc2 (wc2, n_343);
  or g408 (n_424, wc3, n_335);
  not gc3 (wc3, n_336);
  or g409 (n_425, wc4, n_345);
  not gc4 (wc4, n_348);
  or g410 (n_426, wc5, n_390);
  not gc5 (wc5, n_393);
  or g411 (n_427, wc6, n_350);
  not gc6 (wc6, n_353);
  or g412 (n_428, wc7, n_340);
  not gc7 (wc7, n_341);
  or g413 (n_429, wc8, n_355);
  not gc8 (wc8, n_358);
  or g414 (n_430, wc9, n_385);
  not gc9 (wc9, n_388);
  or g415 (n_431, wc10, n_360);
  not gc10 (wc10, n_363);
  or g416 (n_432, wc11, n_365);
  not gc11 (wc11, n_368);
  or g417 (n_433, wc12, n_380);
  not gc12 (wc12, n_383);
  or g418 (n_434, wc13, n_345);
  not gc13 (wc13, n_346);
  or g419 (n_435, wc14, n_370);
  not gc14 (wc14, n_373);
  or g420 (n_436, wc15, n_375);
  not gc15 (wc15, n_378);
  or g421 (n_437, wc16, n_350);
  not gc16 (wc16, n_351);
  or g422 (n_438, wc17, n_355);
  not gc17 (wc17, n_356);
  or g423 (n_439, wc18, n_360);
  not gc18 (wc18, n_361);
  or g424 (n_440, wc19, n_365);
  not gc19 (wc19, n_366);
  or g425 (n_441, wc20, n_370);
  not gc20 (wc20, n_371);
  or g426 (n_442, wc21, n_375);
  not gc21 (wc21, n_376);
  or g427 (n_443, wc22, n_380);
  not gc22 (wc22, n_381);
  or g428 (n_444, wc23, n_385);
  not gc23 (wc23, n_386);
  or g429 (n_445, wc24, n_390);
  not gc24 (wc24, n_391);
endmodule

module mult_unsigned_35_GENERIC(A, B, Z);
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  mult_unsigned_35_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

