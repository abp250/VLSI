library verilog;
use verilog.vl_types.all;
entity ModuleTesting_tb is
end ModuleTesting_tb;
