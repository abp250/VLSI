module csa_tree_add_27_19_group_57_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( in_2 + ( in_0 * in_1 )  )  ;"
  input [7:0] in_0, in_1;
  input [8:0] in_2;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [8:0] in_2;
  wire [16:0] out_0;
  wire n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
  wire n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187;
  wire n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195;
  wire n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203;
  wire n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211;
  wire n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219;
  wire n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227;
  wire n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251;
  wire n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259;
  wire n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267;
  wire n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275;
  wire n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283;
  wire n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291;
  wire n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299;
  wire n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307;
  wire n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315;
  wire n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323;
  wire n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339;
  wire n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347;
  wire n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_389, n_391, n_394, n_396, n_397, n_399, n_401, n_402;
  wire n_404, n_406, n_407, n_409, n_411, n_412, n_414, n_416;
  wire n_417, n_419, n_421, n_422, n_424, n_426, n_427, n_429;
  wire n_431, n_432, n_434, n_436, n_437, n_439, n_441, n_442;
  wire n_444, n_446, n_447, n_449, n_451, n_452, n_454, n_456;
  wire n_457, n_459, n_462, n_465, n_489, n_490, n_492, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  and g1 (n_59, in_0[0], in_1[0]);
  and g2 (n_58, in_0[1], in_1[0]);
  and g3 (n_79, in_0[2], in_1[0]);
  and g4 (n_83, in_0[3], in_1[0]);
  and g5 (n_90, in_0[4], in_1[0]);
  and g6 (n_100, in_0[5], in_1[0]);
  and g7 (n_113, in_0[6], in_1[0]);
  and g8 (n_127, in_0[7], in_1[0]);
  and g9 (n_78, in_0[0], in_1[1]);
  and g10 (n_81, in_0[1], in_1[1]);
  and g11 (n_86, in_0[2], in_1[1]);
  and g12 (n_93, in_0[3], in_1[1]);
  and g13 (n_103, in_0[4], in_1[1]);
  and g14 (n_115, in_0[5], in_1[1]);
  and g15 (n_130, in_0[6], in_1[1]);
  and g16 (n_144, in_0[7], in_1[1]);
  and g17 (n_80, in_0[0], in_1[2]);
  and g18 (n_84, in_0[1], in_1[2]);
  and g19 (n_91, in_0[2], in_1[2]);
  and g20 (n_101, in_0[3], in_1[2]);
  and g21 (n_114, in_0[4], in_1[2]);
  and g22 (n_76, in_0[5], in_1[2]);
  and g23 (n_148, in_0[6], in_1[2]);
  and g24 (n_163, in_0[7], in_1[2]);
  and g25 (n_85, in_0[0], in_1[3]);
  and g26 (n_92, in_0[1], in_1[3]);
  and g27 (n_102, in_0[2], in_1[3]);
  and g28 (n_61, in_0[3], in_1[3]);
  and g29 (n_129, in_0[4], in_1[3]);
  and g30 (n_145, in_0[5], in_1[3]);
  and g31 (n_164, in_0[6], in_1[3]);
  and g32 (n_180, in_0[7], in_1[3]);
  and g33 (n_94, in_0[0], in_1[4]);
  and g34 (n_104, in_0[1], in_1[4]);
  and g35 (n_116, in_0[2], in_1[4]);
  and g36 (n_131, in_0[3], in_1[4]);
  and g37 (n_147, in_0[4], in_1[4]);
  and g38 (n_167, in_0[5], in_1[4]);
  and g39 (n_181, in_0[6], in_1[4]);
  and g40 (n_194, in_0[7], in_1[4]);
  and g41 (n_105, in_0[0], in_1[5]);
  and g42 (n_117, in_0[1], in_1[5]);
  and g43 (n_132, in_0[2], in_1[5]);
  and g44 (n_149, in_0[3], in_1[5]);
  and g45 (n_165, in_0[4], in_1[5]);
  and g46 (n_184, in_0[5], in_1[5]);
  and g47 (n_195, in_0[6], in_1[5]);
  and g48 (n_205, in_0[7], in_1[5]);
  and g49 (n_60, in_0[0], in_1[6]);
  and g50 (n_77, in_0[1], in_1[6]);
  and g51 (n_150, in_0[2], in_1[6]);
  and g52 (n_166, in_0[3], in_1[6]);
  and g53 (n_182, in_0[4], in_1[6]);
  and g54 (n_197, in_0[5], in_1[6]);
  and g55 (n_206, in_0[6], in_1[6]);
  and g56 (n_213, in_0[7], in_1[6]);
  and g57 (n_128, in_0[0], in_1[7]);
  and g58 (n_146, in_0[1], in_1[7]);
  and g59 (n_168, in_0[2], in_1[7]);
  and g60 (n_183, in_0[3], in_1[7]);
  and g61 (n_196, in_0[4], in_1[7]);
  and g62 (n_207, in_0[5], in_1[7]);
  and g63 (n_214, in_0[6], in_1[7]);
  and g64 (n_218, in_0[7], in_1[7]);
  xor g121 (n_75, in_2[1], n_78);
  and g122 (n_57, in_2[1], n_78);
  xor g123 (n_82, in_2[2], n_79);
  and g124 (n_88, in_2[2], n_79);
  xor g125 (n_220, n_80, n_81);
  xor g126 (n_74, n_220, n_82);
  nand g127 (n_221, n_80, n_81);
  nand g128 (n_222, n_82, n_81);
  nand g129 (n_223, n_80, n_82);
  nand g130 (n_56, n_221, n_222, n_223);
  xor g131 (n_87, in_2[3], n_83);
  and g132 (n_96, in_2[3], n_83);
  xor g133 (n_224, n_84, n_85);
  xor g134 (n_89, n_224, n_86);
  nand g135 (n_225, n_84, n_85);
  nand g136 (n_226, n_86, n_85);
  nand g137 (n_227, n_84, n_86);
  nand g138 (n_97, n_225, n_226, n_227);
  xor g139 (n_228, n_87, n_88);
  xor g140 (n_73, n_228, n_89);
  nand g141 (n_229, n_87, n_88);
  nand g142 (n_230, n_89, n_88);
  nand g143 (n_231, n_87, n_89);
  nand g144 (n_55, n_229, n_230, n_231);
  xor g145 (n_95, in_2[4], n_90);
  and g146 (n_106, in_2[4], n_90);
  xor g147 (n_232, n_91, n_92);
  xor g148 (n_98, n_232, n_93);
  nand g149 (n_233, n_91, n_92);
  nand g150 (n_234, n_93, n_92);
  nand g151 (n_235, n_91, n_93);
  nand g152 (n_108, n_233, n_234, n_235);
  xor g153 (n_236, n_94, n_95);
  xor g154 (n_99, n_236, n_96);
  nand g155 (n_237, n_94, n_95);
  nand g156 (n_238, n_96, n_95);
  nand g157 (n_239, n_94, n_96);
  nand g158 (n_110, n_237, n_238, n_239);
  xor g159 (n_240, n_97, n_98);
  xor g160 (n_72, n_240, n_99);
  nand g161 (n_241, n_97, n_98);
  nand g162 (n_242, n_99, n_98);
  nand g163 (n_243, n_97, n_99);
  nand g164 (n_54, n_241, n_242, n_243);
  xor g165 (n_107, in_2[5], n_100);
  and g166 (n_118, in_2[5], n_100);
  xor g167 (n_244, n_101, n_102);
  xor g168 (n_109, n_244, n_103);
  nand g169 (n_245, n_101, n_102);
  nand g170 (n_246, n_103, n_102);
  nand g171 (n_247, n_101, n_103);
  nand g172 (n_120, n_245, n_246, n_247);
  xor g173 (n_248, n_104, n_105);
  xor g174 (n_111, n_248, n_106);
  nand g175 (n_249, n_104, n_105);
  nand g176 (n_250, n_106, n_105);
  nand g177 (n_251, n_104, n_106);
  nand g178 (n_123, n_249, n_250, n_251);
  xor g179 (n_252, n_107, n_108);
  xor g180 (n_112, n_252, n_109);
  nand g181 (n_253, n_107, n_108);
  nand g182 (n_254, n_109, n_108);
  nand g183 (n_255, n_107, n_109);
  nand g184 (n_125, n_253, n_254, n_255);
  xor g185 (n_256, n_110, n_111);
  xor g186 (n_71, n_256, n_112);
  nand g187 (n_257, n_110, n_111);
  nand g188 (n_258, n_112, n_111);
  nand g189 (n_259, n_110, n_112);
  nand g190 (n_53, n_257, n_258, n_259);
  xor g191 (n_119, in_2[6], n_113);
  and g192 (n_134, in_2[6], n_113);
  xor g193 (n_260, n_114, n_60);
  xor g194 (n_122, n_260, n_61);
  nand g195 (n_261, n_114, n_60);
  nand g196 (n_262, n_61, n_60);
  nand g197 (n_263, n_114, n_61);
  nand g198 (n_136, n_261, n_262, n_263);
  xor g199 (n_264, n_115, n_116);
  xor g200 (n_121, n_264, n_117);
  nand g201 (n_265, n_115, n_116);
  nand g202 (n_266, n_117, n_116);
  nand g203 (n_267, n_115, n_117);
  nand g204 (n_135, n_265, n_266, n_267);
  xor g205 (n_268, n_118, n_119);
  xor g206 (n_124, n_268, n_120);
  nand g207 (n_269, n_118, n_119);
  nand g208 (n_270, n_120, n_119);
  nand g209 (n_271, n_118, n_120);
  nand g210 (n_139, n_269, n_270, n_271);
  xor g211 (n_272, n_121, n_122);
  xor g212 (n_126, n_272, n_123);
  nand g213 (n_273, n_121, n_122);
  nand g214 (n_274, n_123, n_122);
  nand g215 (n_275, n_121, n_123);
  nand g216 (n_142, n_273, n_274, n_275);
  xor g217 (n_276, n_124, n_125);
  xor g218 (n_70, n_276, n_126);
  nand g219 (n_277, n_124, n_125);
  nand g220 (n_278, n_126, n_125);
  nand g221 (n_279, n_124, n_126);
  nand g222 (n_52, n_277, n_278, n_279);
  xor g223 (n_133, in_2[7], n_127);
  and g224 (n_151, in_2[7], n_127);
  xor g225 (n_280, n_76, n_77);
  xor g226 (n_138, n_280, n_128);
  nand g227 (n_281, n_76, n_77);
  nand g228 (n_282, n_128, n_77);
  nand g229 (n_283, n_76, n_128);
  nand g230 (n_153, n_281, n_282, n_283);
  xor g231 (n_284, n_129, n_130);
  xor g232 (n_137, n_284, n_131);
  nand g233 (n_285, n_129, n_130);
  nand g234 (n_286, n_131, n_130);
  nand g235 (n_287, n_129, n_131);
  nand g236 (n_154, n_285, n_286, n_287);
  xor g237 (n_288, n_132, n_133);
  xor g238 (n_140, n_288, n_134);
  nand g239 (n_289, n_132, n_133);
  nand g240 (n_290, n_134, n_133);
  nand g241 (n_291, n_132, n_134);
  nand g242 (n_157, n_289, n_290, n_291);
  xor g243 (n_292, n_135, n_136);
  xor g244 (n_141, n_292, n_137);
  nand g245 (n_293, n_135, n_136);
  nand g246 (n_294, n_137, n_136);
  nand g247 (n_295, n_135, n_137);
  nand g248 (n_159, n_293, n_294, n_295);
  xor g249 (n_296, n_138, n_139);
  xor g250 (n_143, n_296, n_140);
  nand g251 (n_297, n_138, n_139);
  nand g252 (n_298, n_140, n_139);
  nand g253 (n_299, n_138, n_140);
  nand g254 (n_161, n_297, n_298, n_299);
  xor g255 (n_300, n_141, n_142);
  xor g256 (n_69, n_300, n_143);
  nand g257 (n_301, n_141, n_142);
  nand g258 (n_302, n_143, n_142);
  nand g259 (n_303, n_141, n_143);
  nand g260 (n_51, n_301, n_302, n_303);
  xor g261 (n_152, in_2[8], n_144);
  and g262 (n_170, in_2[8], n_144);
  xor g263 (n_304, n_145, n_146);
  xor g264 (n_156, n_304, n_147);
  nand g265 (n_305, n_145, n_146);
  nand g266 (n_306, n_147, n_146);
  nand g267 (n_307, n_145, n_147);
  nand g268 (n_171, n_305, n_306, n_307);
  xor g269 (n_308, n_148, n_149);
  xor g270 (n_155, n_308, n_150);
  nand g271 (n_309, n_148, n_149);
  nand g272 (n_310, n_150, n_149);
  nand g273 (n_311, n_148, n_150);
  nand g274 (n_172, n_309, n_310, n_311);
  xor g275 (n_312, n_151, n_152);
  xor g276 (n_158, n_312, n_153);
  nand g277 (n_313, n_151, n_152);
  nand g278 (n_314, n_153, n_152);
  nand g279 (n_315, n_151, n_153);
  nand g280 (n_175, n_313, n_314, n_315);
  xor g281 (n_316, n_154, n_155);
  xor g282 (n_160, n_316, n_156);
  nand g283 (n_317, n_154, n_155);
  nand g284 (n_318, n_156, n_155);
  nand g285 (n_319, n_154, n_156);
  nand g286 (n_176, n_317, n_318, n_319);
  xor g287 (n_320, n_157, n_158);
  xor g288 (n_162, n_320, n_159);
  nand g289 (n_321, n_157, n_158);
  nand g290 (n_322, n_159, n_158);
  nand g291 (n_323, n_157, n_159);
  nand g292 (n_179, n_321, n_322, n_323);
  xor g293 (n_324, n_160, n_161);
  xor g294 (n_68, n_324, n_162);
  nand g295 (n_325, n_160, n_161);
  nand g296 (n_326, n_162, n_161);
  nand g297 (n_327, n_160, n_162);
  nand g298 (n_50, n_325, n_326, n_327);
  xor g299 (n_169, n_163, n_164);
  and g300 (n_186, n_163, n_164);
  xor g301 (n_328, n_165, n_166);
  xor g302 (n_173, n_328, n_167);
  nand g303 (n_329, n_165, n_166);
  nand g304 (n_330, n_167, n_166);
  nand g305 (n_331, n_165, n_167);
  nand g306 (n_187, n_329, n_330, n_331);
  xor g307 (n_332, n_168, n_169);
  xor g308 (n_174, n_332, n_170);
  nand g309 (n_333, n_168, n_169);
  nand g310 (n_334, n_170, n_169);
  nand g311 (n_335, n_168, n_170);
  nand g312 (n_189, n_333, n_334, n_335);
  xor g313 (n_336, n_171, n_172);
  xor g314 (n_177, n_336, n_173);
  nand g315 (n_337, n_171, n_172);
  nand g316 (n_338, n_173, n_172);
  nand g317 (n_339, n_171, n_173);
  nand g318 (n_191, n_337, n_338, n_339);
  xor g319 (n_340, n_174, n_175);
  xor g320 (n_178, n_340, n_176);
  nand g321 (n_341, n_174, n_175);
  nand g322 (n_342, n_176, n_175);
  nand g323 (n_343, n_174, n_176);
  nand g324 (n_193, n_341, n_342, n_343);
  xor g325 (n_344, n_177, n_178);
  xor g326 (n_67, n_344, n_179);
  nand g327 (n_345, n_177, n_178);
  nand g328 (n_346, n_179, n_178);
  nand g329 (n_347, n_177, n_179);
  nand g330 (n_49, n_345, n_346, n_347);
  xor g331 (n_185, n_180, n_181);
  and g332 (n_198, n_180, n_181);
  xor g333 (n_348, n_182, n_183);
  xor g334 (n_188, n_348, n_184);
  nand g335 (n_349, n_182, n_183);
  nand g336 (n_350, n_184, n_183);
  nand g337 (n_351, n_182, n_184);
  nand g338 (n_200, n_349, n_350, n_351);
  xor g339 (n_352, n_185, n_186);
  xor g340 (n_190, n_352, n_187);
  nand g341 (n_353, n_185, n_186);
  nand g342 (n_354, n_187, n_186);
  nand g343 (n_355, n_185, n_187);
  nand g344 (n_202, n_353, n_354, n_355);
  xor g345 (n_356, n_188, n_189);
  xor g346 (n_192, n_356, n_190);
  nand g347 (n_357, n_188, n_189);
  nand g348 (n_358, n_190, n_189);
  nand g349 (n_359, n_188, n_190);
  nand g350 (n_204, n_357, n_358, n_359);
  xor g351 (n_360, n_191, n_192);
  xor g352 (n_66, n_360, n_193);
  nand g353 (n_361, n_191, n_192);
  nand g354 (n_362, n_193, n_192);
  nand g355 (n_363, n_191, n_193);
  nand g356 (n_65, n_361, n_362, n_363);
  xor g357 (n_199, n_194, n_195);
  and g358 (n_208, n_194, n_195);
  xor g359 (n_364, n_196, n_197);
  xor g360 (n_201, n_364, n_198);
  nand g361 (n_365, n_196, n_197);
  nand g362 (n_366, n_198, n_197);
  nand g363 (n_367, n_196, n_198);
  nand g364 (n_210, n_365, n_366, n_367);
  xor g365 (n_368, n_199, n_200);
  xor g366 (n_203, n_368, n_201);
  nand g367 (n_369, n_199, n_200);
  nand g368 (n_370, n_201, n_200);
  nand g369 (n_371, n_199, n_201);
  nand g370 (n_212, n_369, n_370, n_371);
  xor g371 (n_372, n_202, n_203);
  xor g372 (n_48, n_372, n_204);
  nand g373 (n_373, n_202, n_203);
  nand g374 (n_374, n_204, n_203);
  nand g375 (n_375, n_202, n_204);
  nand g376 (n_64, n_373, n_374, n_375);
  xor g377 (n_209, n_205, n_206);
  and g378 (n_215, n_205, n_206);
  xor g379 (n_376, n_207, n_208);
  xor g380 (n_211, n_376, n_209);
  nand g381 (n_377, n_207, n_208);
  nand g382 (n_378, n_209, n_208);
  nand g383 (n_379, n_207, n_209);
  nand g384 (n_217, n_377, n_378, n_379);
  xor g385 (n_380, n_210, n_211);
  xor g386 (n_47, n_380, n_212);
  nand g387 (n_381, n_210, n_211);
  nand g388 (n_382, n_212, n_211);
  nand g389 (n_383, n_210, n_212);
  nand g390 (n_63, n_381, n_382, n_383);
  xor g391 (n_216, n_213, n_214);
  and g392 (n_219, n_213, n_214);
  xor g393 (n_384, n_215, n_216);
  xor g394 (n_46, n_384, n_217);
  nand g395 (n_385, n_215, n_216);
  nand g396 (n_386, n_217, n_216);
  nand g397 (n_387, n_215, n_217);
  nand g398 (n_62, n_385, n_386, n_387);
  xor g399 (n_45, n_218, n_219);
  and g400 (n_44, n_218, n_219);
  nand g403 (n_389, n_59, in_2[0]);
  nor g406 (n_391, n_58, n_75);
  nand g407 (n_394, n_58, n_75);
  nor g408 (n_396, n_57, n_74);
  nand g409 (n_399, n_57, n_74);
  nor g410 (n_401, n_56, n_73);
  nand g411 (n_404, n_56, n_73);
  nor g412 (n_406, n_55, n_72);
  nand g413 (n_409, n_55, n_72);
  nor g414 (n_411, n_54, n_71);
  nand g415 (n_414, n_54, n_71);
  nor g416 (n_416, n_53, n_70);
  nand g417 (n_419, n_53, n_70);
  nor g418 (n_421, n_52, n_69);
  nand g419 (n_424, n_52, n_69);
  nor g420 (n_426, n_51, n_68);
  nand g421 (n_429, n_51, n_68);
  nor g422 (n_431, n_50, n_67);
  nand g423 (n_434, n_50, n_67);
  nor g424 (n_436, n_49, n_66);
  nand g425 (n_439, n_49, n_66);
  nor g426 (n_441, n_48, n_65);
  nand g427 (n_444, n_48, n_65);
  nor g428 (n_446, n_47, n_64);
  nand g429 (n_449, n_47, n_64);
  nor g430 (n_451, n_46, n_63);
  nand g431 (n_454, n_46, n_63);
  nor g432 (n_456, n_45, n_62);
  nand g433 (n_459, n_45, n_62);
  nand g440 (n_397, n_394, n_489);
  nand g443 (n_402, n_399, n_494);
  nand g446 (n_407, n_404, n_497);
  nand g449 (n_412, n_409, n_502);
  nand g452 (n_417, n_414, n_509);
  nand g455 (n_422, n_419, n_510);
  nand g458 (n_427, n_424, n_511);
  nand g461 (n_432, n_429, n_512);
  nand g464 (n_437, n_434, n_513);
  nand g67 (n_442, n_439, n_514);
  nand g70 (n_447, n_444, n_515);
  nand g73 (n_452, n_449, n_516);
  nand g76 (n_457, n_454, n_517);
  nand g79 (n_462, n_459, n_518);
  nand g81 (n_465, n_462, n_44);
  xnor g89 (out_0[2], n_397, n_492);
  xnor g91 (out_0[3], n_402, n_495);
  xnor g93 (out_0[4], n_407, n_496);
  xnor g95 (out_0[5], n_412, n_498);
  xnor g97 (out_0[6], n_417, n_500);
  xnor g99 (out_0[7], n_422, n_503);
  xnor g101 (out_0[8], n_427, n_505);
  xnor g103 (out_0[9], n_432, n_506);
  xnor g105 (out_0[10], n_437, n_507);
  xnor g107 (out_0[11], n_442, n_508);
  xnor g109 (out_0[12], n_447, n_504);
  xnor g111 (out_0[13], n_452, n_501);
  xnor g113 (out_0[14], n_457, n_499);
  xor g118 (out_0[0], in_2[0], n_59);
  or g467 (n_489, n_389, n_391);
  or g468 (n_490, wc, n_391);
  not gc (wc, n_394);
  xor g469 (out_0[1], n_389, n_490);
  or g470 (n_492, wc0, n_396);
  not gc0 (wc0, n_399);
  or g472 (n_494, wc1, n_396);
  not gc1 (wc1, n_397);
  or g473 (n_495, wc2, n_401);
  not gc2 (wc2, n_404);
  or g474 (n_496, wc3, n_406);
  not gc3 (wc3, n_409);
  or g475 (n_497, wc4, n_401);
  not gc4 (wc4, n_402);
  or g476 (n_498, wc5, n_411);
  not gc5 (wc5, n_414);
  or g477 (n_499, wc6, n_456);
  not gc6 (wc6, n_459);
  or g478 (n_500, wc7, n_416);
  not gc7 (wc7, n_419);
  or g479 (n_501, wc8, n_451);
  not gc8 (wc8, n_454);
  or g480 (n_502, wc9, n_406);
  not gc9 (wc9, n_407);
  or g481 (n_503, wc10, n_421);
  not gc10 (wc10, n_424);
  or g482 (n_504, wc11, n_446);
  not gc11 (wc11, n_449);
  or g483 (n_505, wc12, n_426);
  not gc12 (wc12, n_429);
  or g484 (n_506, wc13, n_431);
  not gc13 (wc13, n_434);
  or g485 (n_507, wc14, n_436);
  not gc14 (wc14, n_439);
  or g486 (n_508, wc15, n_441);
  not gc15 (wc15, n_444);
  or g487 (n_509, wc16, n_411);
  not gc16 (wc16, n_412);
  or g488 (n_510, wc17, n_416);
  not gc17 (wc17, n_417);
  or g489 (n_511, wc18, n_421);
  not gc18 (wc18, n_422);
  or g490 (n_512, wc19, n_426);
  not gc19 (wc19, n_427);
  or g491 (n_513, wc20, n_431);
  not gc20 (wc20, n_432);
  or g492 (n_514, wc21, n_436);
  not gc21 (wc21, n_437);
  or g493 (n_515, wc22, n_441);
  not gc22 (wc22, n_442);
  or g494 (n_516, wc23, n_446);
  not gc23 (wc23, n_447);
  or g495 (n_517, wc24, n_451);
  not gc24 (wc24, n_452);
  or g496 (n_518, wc25, n_456);
  not gc25 (wc25, n_457);
  xor g497 (out_0[15], n_44, n_462);
  not g498 (out_0[16], n_465);
endmodule

module csa_tree_add_27_19_group_57_GENERIC(in_0, in_1, in_2, out_0);
  input [7:0] in_0, in_1;
  input [8:0] in_2;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [8:0] in_2;
  wire [16:0] out_0;
  csa_tree_add_27_19_group_57_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module mult_unsigned_85_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $unsigned(A) * $unsigned(B);"
  input [7:0] A, B;
  output [7:0] Z;
  wire [7:0] A, B;
  wire [7:0] Z;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_33;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_142, n_146, n_150, n_154, n_161, n_164, n_166, n_169;
  wire n_171, n_172, n_174, n_176, n_177, n_179, n_181, n_182;
  wire n_184, n_186, n_187, n_189, n_191, n_192, n_194, n_206;
  wire n_208, n_209, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219;
  and g1 (Z[0], A[0], B[0]);
  and g2 (n_31, A[1], B[0]);
  and g3 (n_42, A[2], B[0]);
  and g4 (n_44, A[3], B[0]);
  and g5 (n_49, A[4], B[0]);
  and g6 (n_41, A[5], B[0]);
  and g7 (n_67, A[6], B[0]);
  and g8 (n_81, A[7], B[0]);
  and g9 (n_39, A[0], B[1]);
  and g10 (n_30, A[1], B[1]);
  and g11 (n_45, A[2], B[1]);
  and g12 (n_50, A[3], B[1]);
  and g13 (n_57, A[4], B[1]);
  and g14 (n_68, A[5], B[1]);
  and g15 (n_82, A[6], B[1]);
  and g16 (n_43, A[0], B[2]);
  and g17 (n_47, A[1], B[2]);
  and g18 (n_53, A[2], B[2]);
  and g19 (n_60, A[3], B[2]);
  and g20 (n_71, A[4], B[2]);
  and g21 (n_86, A[5], B[2]);
  and g22 (n_46, A[0], B[3]);
  and g23 (n_51, A[1], B[3]);
  and g24 (n_58, A[2], B[3]);
  and g25 (n_69, A[3], B[3]);
  and g26 (n_83, A[4], B[3]);
  and g27 (n_52, A[0], B[4]);
  and g28 (n_59, A[1], B[4]);
  and g29 (n_70, A[2], B[4]);
  and g30 (n_85, A[3], B[4]);
  and g31 (n_61, A[0], B[5]);
  and g32 (n_72, A[1], B[5]);
  and g33 (n_87, A[2], B[5]);
  and g34 (n_73, A[0], B[6]);
  and g35 (n_88, A[1], B[6]);
  and g36 (n_84, A[0], B[7]);
  xor g58 (n_38, n_42, n_43);
  and g59 (n_29, n_42, n_43);
  xor g60 (n_48, n_44, n_45);
  and g61 (n_55, n_44, n_45);
  xor g62 (n_98, n_46, n_47);
  xor g63 (n_37, n_98, n_48);
  nand g64 (n_99, n_46, n_47);
  nand g65 (n_100, n_48, n_47);
  nand g66 (n_101, n_46, n_48);
  nand g67 (n_28, n_99, n_100, n_101);
  xor g68 (n_54, n_49, n_50);
  and g69 (n_63, n_49, n_50);
  xor g70 (n_102, n_51, n_52);
  xor g71 (n_56, n_102, n_53);
  nand g72 (n_103, n_51, n_52);
  nand g73 (n_104, n_53, n_52);
  nand g74 (n_105, n_51, n_53);
  nand g75 (n_64, n_103, n_104, n_105);
  xor g76 (n_106, n_54, n_55);
  xor g77 (n_36, n_106, n_56);
  nand g78 (n_107, n_54, n_55);
  nand g79 (n_108, n_56, n_55);
  nand g80 (n_109, n_54, n_56);
  nand g81 (n_27, n_107, n_108, n_109);
  xor g82 (n_62, n_41, n_57);
  and g83 (n_74, n_41, n_57);
  xor g84 (n_110, n_58, n_59);
  xor g85 (n_65, n_110, n_60);
  nand g86 (n_111, n_58, n_59);
  nand g87 (n_112, n_60, n_59);
  nand g88 (n_113, n_58, n_60);
  nand g89 (n_76, n_111, n_112, n_113);
  xor g90 (n_114, n_61, n_62);
  xor g91 (n_66, n_114, n_63);
  nand g92 (n_115, n_61, n_62);
  nand g93 (n_116, n_63, n_62);
  nand g94 (n_117, n_61, n_63);
  nand g95 (n_78, n_115, n_116, n_117);
  xor g96 (n_118, n_64, n_65);
  xor g97 (n_35, n_118, n_66);
  nand g98 (n_119, n_64, n_65);
  nand g99 (n_120, n_66, n_65);
  nand g100 (n_121, n_64, n_66);
  nand g101 (n_26, n_119, n_120, n_121);
  xor g102 (n_75, n_67, n_68);
  and g103 (n_89, n_67, n_68);
  xor g104 (n_122, n_69, n_70);
  xor g105 (n_77, n_122, n_71);
  nand g106 (n_123, n_69, n_70);
  nand g107 (n_124, n_71, n_70);
  nand g108 (n_125, n_69, n_71);
  nand g109 (n_91, n_123, n_124, n_125);
  xor g110 (n_126, n_72, n_73);
  xor g111 (n_79, n_126, n_74);
  nand g112 (n_127, n_72, n_73);
  nand g113 (n_128, n_74, n_73);
  nand g114 (n_129, n_72, n_74);
  nand g115 (n_94, n_127, n_128, n_129);
  xor g116 (n_130, n_75, n_76);
  xor g117 (n_80, n_130, n_77);
  nand g118 (n_131, n_75, n_76);
  nand g119 (n_132, n_77, n_76);
  nand g120 (n_133, n_75, n_77);
  nand g121 (n_96, n_131, n_132, n_133);
  xor g122 (n_134, n_78, n_79);
  xor g123 (n_34, n_134, n_80);
  nand g124 (n_135, n_78, n_79);
  nand g125 (n_136, n_80, n_79);
  nand g126 (n_137, n_78, n_80);
  nand g127 (n_25, n_135, n_136, n_137);
  xor g128 (n_90, n_81, n_82);
  xor g130 (n_138, n_83, n_84);
  xor g131 (n_93, n_138, n_85);
  xor g136 (n_142, n_86, n_87);
  xor g137 (n_92, n_142, n_88);
  xor g142 (n_146, n_89, n_90);
  xor g143 (n_95, n_146, n_91);
  xor g148 (n_150, n_92, n_93);
  xor g149 (n_97, n_150, n_94);
  xor g154 (n_154, n_95, n_96);
  xor g155 (n_33, n_154, n_97);
  nor g165 (n_161, n_31, n_39);
  nand g166 (n_164, n_31, n_39);
  nor g167 (n_166, n_30, n_38);
  nand g168 (n_169, n_30, n_38);
  nor g169 (n_171, n_29, n_37);
  nand g170 (n_174, n_29, n_37);
  nor g171 (n_176, n_28, n_36);
  nand g172 (n_179, n_28, n_36);
  nor g173 (n_181, n_27, n_35);
  nand g174 (n_184, n_27, n_35);
  nor g175 (n_186, n_26, n_34);
  nand g176 (n_189, n_26, n_34);
  nor g177 (n_191, n_25, n_33);
  nand g178 (n_194, n_25, n_33);
  nand g184 (n_172, n_169, n_209);
  nand g187 (n_177, n_174, n_213);
  nand g190 (n_182, n_179, n_216);
  nand g193 (n_187, n_184, n_218);
  nand g37 (n_192, n_189, n_219);
  xnor g46 (Z[3], n_172, n_211);
  xnor g48 (Z[4], n_177, n_212);
  xnor g50 (Z[5], n_182, n_214);
  xnor g52 (Z[6], n_187, n_215);
  xnor g54 (Z[7], n_192, n_217);
  or g196 (n_206, wc, n_161);
  not gc (wc, n_164);
  not g198 (Z[1], n_206);
  or g199 (n_208, wc0, n_166);
  not gc0 (wc0, n_169);
  or g200 (n_209, n_164, n_166);
  xor g201 (Z[2], n_164, n_208);
  or g202 (n_211, wc1, n_171);
  not gc1 (wc1, n_174);
  or g203 (n_212, wc2, n_176);
  not gc2 (wc2, n_179);
  or g204 (n_213, wc3, n_171);
  not gc3 (wc3, n_172);
  or g205 (n_214, wc4, n_181);
  not gc4 (wc4, n_184);
  or g206 (n_215, wc5, n_186);
  not gc5 (wc5, n_189);
  or g207 (n_216, wc6, n_176);
  not gc6 (wc6, n_177);
  or g208 (n_217, wc7, n_191);
  not gc7 (wc7, n_194);
  or g209 (n_218, wc8, n_181);
  not gc8 (wc8, n_182);
  or g210 (n_219, wc9, n_186);
  not gc9 (wc9, n_187);
endmodule

module mult_unsigned_85_GENERIC(A, B, Z);
  input [7:0] A, B;
  output [7:0] Z;
  wire [7:0] A, B;
  wire [7:0] Z;
  mult_unsigned_85_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

