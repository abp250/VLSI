module add_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [15:0] A, B;
  output [15:0] Z;
  wire [15:0] A, B;
  wire [15:0] Z;
  wire n_50, n_53, n_56, n_58, n_59, n_60, n_61, n_63;
  wire n_64, n_65, n_66, n_67, n_69, n_70, n_71, n_72;
  wire n_73, n_75, n_76, n_77, n_78, n_79, n_81, n_82;
  wire n_83, n_84, n_85, n_87, n_88, n_89, n_90, n_91;
  wire n_93, n_94, n_95, n_96, n_99, n_100, n_103, n_105;
  wire n_106, n_107, n_109, n_111, n_116, n_117, n_119, n_121;
  wire n_126, n_127, n_129, n_136, n_139, n_144, n_148, n_149;
  wire n_151, n_155, n_157, n_163, n_166, n_173, n_175, n_178;
  wire n_179, n_181, n_188, n_192, n_194, n_197, n_201, n_203;
  wire n_206, n_209, n_212, n_214, n_217, n_225, n_226, n_227;
  wire n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_245, n_246, n_247, n_248, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_50, A[0], B[0]);
  nor g6 (n_53, A[1], B[1]);
  nand g7 (n_56, A[1], B[1]);
  nor g8 (n_63, A[2], B[2]);
  nand g9 (n_58, A[2], B[2]);
  nor g10 (n_59, A[3], B[3]);
  nand g11 (n_60, A[3], B[3]);
  nor g12 (n_69, A[4], B[4]);
  nand g13 (n_64, A[4], B[4]);
  nor g14 (n_65, A[5], B[5]);
  nand g15 (n_66, A[5], B[5]);
  nor g16 (n_75, A[6], B[6]);
  nand g17 (n_70, A[6], B[6]);
  nor g18 (n_71, A[7], B[7]);
  nand g19 (n_72, A[7], B[7]);
  nor g20 (n_81, A[8], B[8]);
  nand g21 (n_76, A[8], B[8]);
  nor g22 (n_77, A[9], B[9]);
  nand g23 (n_78, A[9], B[9]);
  nor g24 (n_87, A[10], B[10]);
  nand g25 (n_82, A[10], B[10]);
  nor g26 (n_83, A[11], B[11]);
  nand g27 (n_84, A[11], B[11]);
  nor g28 (n_93, A[12], B[12]);
  nand g29 (n_88, A[12], B[12]);
  nor g30 (n_89, A[13], B[13]);
  nand g31 (n_90, A[13], B[13]);
  nor g32 (n_99, A[14], B[14]);
  nand g33 (n_94, A[14], B[14]);
  nor g34 (n_95, A[15], B[15]);
  nand g35 (n_96, A[15], B[15]);
  nand g38 (n_100, n_56, n_225);
  nor g39 (n_61, n_58, n_59);
  nor g42 (n_103, n_63, n_59);
  nor g43 (n_67, n_64, n_65);
  nor g46 (n_109, n_69, n_65);
  nor g47 (n_73, n_70, n_71);
  nor g50 (n_111, n_75, n_71);
  nor g51 (n_79, n_76, n_77);
  nor g54 (n_119, n_81, n_77);
  nor g55 (n_85, n_82, n_83);
  nor g58 (n_121, n_87, n_83);
  nor g59 (n_91, n_88, n_89);
  nor g62 (n_129, n_93, n_89);
  nand g69 (n_188, n_58, n_250);
  nand g70 (n_105, n_103, n_100);
  nand g71 (n_136, n_226, n_105);
  nor g72 (n_107, n_75, n_106);
  nand g81 (n_144, n_109, n_111);
  nor g82 (n_117, n_87, n_116);
  nand g91 (n_151, n_119, n_121);
  nor g92 (n_127, n_99, n_126);
  nand g104 (n_192, n_64, n_256);
  nand g105 (n_139, n_109, n_136);
  nand g106 (n_194, n_106, n_139);
  nand g109 (n_197, n_251, n_257);
  nand g112 (n_163, n_252, n_258);
  nor g113 (n_149, n_93, n_148);
  nor g116 (n_173, n_93, n_151);
  nor g122 (n_157, n_155, n_148);
  nor g125 (n_179, n_151, n_155);
  nand g132 (n_201, n_76, n_262);
  nand g133 (n_166, n_119, n_163);
  nand g134 (n_203, n_116, n_166);
  nand g137 (n_206, n_253, n_263);
  nand g140 (n_209, n_148, n_264);
  nand g141 (n_175, n_173, n_163);
  nand g142 (n_212, n_259, n_175);
  nand g143 (n_178, n_248, n_163);
  nand g144 (n_214, n_260, n_178);
  nand g145 (n_181, n_179, n_163);
  nand g146 (n_217, n_261, n_181);
  xnor g152 (Z[2], n_100, n_232);
  xnor g155 (Z[3], n_188, n_233);
  xnor g157 (Z[4], n_136, n_234);
  xnor g160 (Z[5], n_192, n_235);
  xnor g162 (Z[6], n_194, n_236);
  xnor g165 (Z[7], n_197, n_237);
  xnor g167 (Z[8], n_163, n_238);
  xnor g170 (Z[9], n_201, n_239);
  xnor g172 (Z[10], n_203, n_240);
  xnor g175 (Z[11], n_206, n_241);
  xnor g178 (Z[12], n_209, n_242);
  xnor g181 (Z[13], n_212, n_243);
  xnor g183 (Z[14], n_214, n_244);
  xnor g186 (Z[15], n_217, n_245);
  or g189 (n_225, n_50, n_53);
  and g190 (n_226, wc, n_60);
  not gc (wc, n_61);
  and g191 (n_106, wc0, n_66);
  not gc0 (wc0, n_67);
  and g192 (n_227, wc1, n_72);
  not gc1 (wc1, n_73);
  and g193 (n_116, wc2, n_78);
  not gc2 (wc2, n_79);
  and g194 (n_228, wc3, n_84);
  not gc3 (wc3, n_85);
  and g195 (n_126, wc4, n_90);
  not gc4 (wc4, n_91);
  or g196 (n_229, wc5, n_75);
  not gc5 (wc5, n_109);
  or g197 (n_230, wc6, n_87);
  not gc6 (wc6, n_119);
  or g198 (n_155, wc7, n_99);
  not gc7 (wc7, n_129);
  or g199 (n_231, wc8, n_53);
  not gc8 (wc8, n_56);
  or g200 (n_232, wc9, n_63);
  not gc9 (wc9, n_58);
  or g201 (n_233, wc10, n_59);
  not gc10 (wc10, n_60);
  or g202 (n_234, wc11, n_69);
  not gc11 (wc11, n_64);
  or g203 (n_235, wc12, n_65);
  not gc12 (wc12, n_66);
  or g204 (n_236, wc13, n_75);
  not gc13 (wc13, n_70);
  or g205 (n_237, wc14, n_71);
  not gc14 (wc14, n_72);
  or g206 (n_238, wc15, n_81);
  not gc15 (wc15, n_76);
  or g207 (n_239, wc16, n_77);
  not gc16 (wc16, n_78);
  or g208 (n_240, wc17, n_87);
  not gc17 (wc17, n_82);
  or g209 (n_241, wc18, n_83);
  not gc18 (wc18, n_84);
  or g210 (n_242, wc19, n_93);
  not gc19 (wc19, n_88);
  or g211 (n_243, wc20, n_89);
  not gc20 (wc20, n_90);
  or g212 (n_244, wc21, n_99);
  not gc21 (wc21, n_94);
  or g213 (n_245, wc22, n_95);
  not gc22 (wc22, n_96);
  and g214 (n_246, wc23, n_111);
  not gc23 (wc23, n_106);
  and g215 (n_247, wc24, n_121);
  not gc24 (wc24, n_116);
  and g216 (n_248, wc25, n_129);
  not gc25 (wc25, n_151);
  xor g217 (Z[1], n_50, n_231);
  or g218 (n_250, wc26, n_63);
  not gc26 (wc26, n_100);
  and g219 (n_251, wc27, n_70);
  not gc27 (wc27, n_107);
  and g220 (n_252, wc28, n_227);
  not gc28 (wc28, n_246);
  and g221 (n_253, wc29, n_82);
  not gc29 (wc29, n_117);
  and g222 (n_148, wc30, n_228);
  not gc30 (wc30, n_247);
  and g223 (n_254, wc31, n_94);
  not gc31 (wc31, n_127);
  and g224 (n_255, wc32, n_129);
  not gc32 (wc32, n_148);
  or g225 (n_256, wc33, n_69);
  not gc33 (wc33, n_136);
  or g226 (n_257, n_229, wc34);
  not gc34 (wc34, n_136);
  or g227 (n_258, n_144, wc35);
  not gc35 (wc35, n_136);
  and g228 (n_259, wc36, n_88);
  not gc36 (wc36, n_149);
  and g229 (n_260, wc37, n_126);
  not gc37 (wc37, n_255);
  and g230 (n_261, n_254, wc38);
  not gc38 (wc38, n_157);
  or g231 (n_262, wc39, n_81);
  not gc39 (wc39, n_163);
  or g232 (n_263, n_230, wc40);
  not gc40 (wc40, n_163);
  or g233 (n_264, wc41, n_151);
  not gc41 (wc41, n_163);
endmodule

module add_unsigned_GENERIC(A, B, Z);
  input [15:0] A, B;
  output [15:0] Z;
  wire [15:0] A, B;
  wire [15:0] Z;
  add_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_32_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [15:0] A, B;
  output [15:0] Z;
  wire [15:0] A, B;
  wire [15:0] Z;
  wire n_50, n_53, n_56, n_58, n_59, n_60, n_61, n_63;
  wire n_64, n_65, n_66, n_67, n_69, n_70, n_71, n_72;
  wire n_73, n_75, n_76, n_77, n_78, n_79, n_81, n_82;
  wire n_83, n_84, n_85, n_87, n_88, n_89, n_90, n_91;
  wire n_93, n_94, n_95, n_96, n_99, n_100, n_103, n_105;
  wire n_106, n_107, n_109, n_111, n_116, n_117, n_119, n_121;
  wire n_126, n_127, n_129, n_136, n_139, n_144, n_148, n_149;
  wire n_151, n_155, n_157, n_163, n_166, n_173, n_175, n_178;
  wire n_179, n_181, n_188, n_192, n_194, n_197, n_201, n_203;
  wire n_206, n_209, n_212, n_214, n_217, n_225, n_226, n_227;
  wire n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_245, n_246, n_247, n_248, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264;
  xor g1 (Z[0], A[0], B[0]);
  nand g2 (n_50, A[0], B[0]);
  nor g6 (n_53, A[1], B[1]);
  nand g7 (n_56, A[1], B[1]);
  nor g8 (n_63, A[2], B[2]);
  nand g9 (n_58, A[2], B[2]);
  nor g10 (n_59, A[3], B[3]);
  nand g11 (n_60, A[3], B[3]);
  nor g12 (n_69, A[4], B[4]);
  nand g13 (n_64, A[4], B[4]);
  nor g14 (n_65, A[5], B[5]);
  nand g15 (n_66, A[5], B[5]);
  nor g16 (n_75, A[6], B[6]);
  nand g17 (n_70, A[6], B[6]);
  nor g18 (n_71, A[7], B[7]);
  nand g19 (n_72, A[7], B[7]);
  nor g20 (n_81, A[8], B[8]);
  nand g21 (n_76, A[8], B[8]);
  nor g22 (n_77, A[9], B[9]);
  nand g23 (n_78, A[9], B[9]);
  nor g24 (n_87, A[10], B[10]);
  nand g25 (n_82, A[10], B[10]);
  nor g26 (n_83, A[11], B[11]);
  nand g27 (n_84, A[11], B[11]);
  nor g28 (n_93, A[12], B[12]);
  nand g29 (n_88, A[12], B[12]);
  nor g30 (n_89, A[13], B[13]);
  nand g31 (n_90, A[13], B[13]);
  nor g32 (n_99, A[14], B[14]);
  nand g33 (n_94, A[14], B[14]);
  nor g34 (n_95, A[15], B[15]);
  nand g35 (n_96, A[15], B[15]);
  nand g38 (n_100, n_56, n_225);
  nor g39 (n_61, n_58, n_59);
  nor g42 (n_103, n_63, n_59);
  nor g43 (n_67, n_64, n_65);
  nor g46 (n_109, n_69, n_65);
  nor g47 (n_73, n_70, n_71);
  nor g50 (n_111, n_75, n_71);
  nor g51 (n_79, n_76, n_77);
  nor g54 (n_119, n_81, n_77);
  nor g55 (n_85, n_82, n_83);
  nor g58 (n_121, n_87, n_83);
  nor g59 (n_91, n_88, n_89);
  nor g62 (n_129, n_93, n_89);
  nand g69 (n_188, n_58, n_250);
  nand g70 (n_105, n_103, n_100);
  nand g71 (n_136, n_226, n_105);
  nor g72 (n_107, n_75, n_106);
  nand g81 (n_144, n_109, n_111);
  nor g82 (n_117, n_87, n_116);
  nand g91 (n_151, n_119, n_121);
  nor g92 (n_127, n_99, n_126);
  nand g104 (n_192, n_64, n_256);
  nand g105 (n_139, n_109, n_136);
  nand g106 (n_194, n_106, n_139);
  nand g109 (n_197, n_251, n_257);
  nand g112 (n_163, n_252, n_258);
  nor g113 (n_149, n_93, n_148);
  nor g116 (n_173, n_93, n_151);
  nor g122 (n_157, n_155, n_148);
  nor g125 (n_179, n_151, n_155);
  nand g132 (n_201, n_76, n_262);
  nand g133 (n_166, n_119, n_163);
  nand g134 (n_203, n_116, n_166);
  nand g137 (n_206, n_253, n_263);
  nand g140 (n_209, n_148, n_264);
  nand g141 (n_175, n_173, n_163);
  nand g142 (n_212, n_259, n_175);
  nand g143 (n_178, n_248, n_163);
  nand g144 (n_214, n_260, n_178);
  nand g145 (n_181, n_179, n_163);
  nand g146 (n_217, n_261, n_181);
  xnor g152 (Z[2], n_100, n_232);
  xnor g155 (Z[3], n_188, n_233);
  xnor g157 (Z[4], n_136, n_234);
  xnor g160 (Z[5], n_192, n_235);
  xnor g162 (Z[6], n_194, n_236);
  xnor g165 (Z[7], n_197, n_237);
  xnor g167 (Z[8], n_163, n_238);
  xnor g170 (Z[9], n_201, n_239);
  xnor g172 (Z[10], n_203, n_240);
  xnor g175 (Z[11], n_206, n_241);
  xnor g178 (Z[12], n_209, n_242);
  xnor g181 (Z[13], n_212, n_243);
  xnor g183 (Z[14], n_214, n_244);
  xnor g186 (Z[15], n_217, n_245);
  or g189 (n_225, n_50, n_53);
  and g190 (n_226, wc, n_60);
  not gc (wc, n_61);
  and g191 (n_106, wc0, n_66);
  not gc0 (wc0, n_67);
  and g192 (n_227, wc1, n_72);
  not gc1 (wc1, n_73);
  and g193 (n_116, wc2, n_78);
  not gc2 (wc2, n_79);
  and g194 (n_228, wc3, n_84);
  not gc3 (wc3, n_85);
  and g195 (n_126, wc4, n_90);
  not gc4 (wc4, n_91);
  or g196 (n_229, wc5, n_75);
  not gc5 (wc5, n_109);
  or g197 (n_230, wc6, n_87);
  not gc6 (wc6, n_119);
  or g198 (n_155, wc7, n_99);
  not gc7 (wc7, n_129);
  or g199 (n_231, wc8, n_53);
  not gc8 (wc8, n_56);
  or g200 (n_232, wc9, n_63);
  not gc9 (wc9, n_58);
  or g201 (n_233, wc10, n_59);
  not gc10 (wc10, n_60);
  or g202 (n_234, wc11, n_69);
  not gc11 (wc11, n_64);
  or g203 (n_235, wc12, n_65);
  not gc12 (wc12, n_66);
  or g204 (n_236, wc13, n_75);
  not gc13 (wc13, n_70);
  or g205 (n_237, wc14, n_71);
  not gc14 (wc14, n_72);
  or g206 (n_238, wc15, n_81);
  not gc15 (wc15, n_76);
  or g207 (n_239, wc16, n_77);
  not gc16 (wc16, n_78);
  or g208 (n_240, wc17, n_87);
  not gc17 (wc17, n_82);
  or g209 (n_241, wc18, n_83);
  not gc18 (wc18, n_84);
  or g210 (n_242, wc19, n_93);
  not gc19 (wc19, n_88);
  or g211 (n_243, wc20, n_89);
  not gc20 (wc20, n_90);
  or g212 (n_244, wc21, n_99);
  not gc21 (wc21, n_94);
  or g213 (n_245, wc22, n_95);
  not gc22 (wc22, n_96);
  and g214 (n_246, wc23, n_111);
  not gc23 (wc23, n_106);
  and g215 (n_247, wc24, n_121);
  not gc24 (wc24, n_116);
  and g216 (n_248, wc25, n_129);
  not gc25 (wc25, n_151);
  xor g217 (Z[1], n_50, n_231);
  or g218 (n_250, wc26, n_63);
  not gc26 (wc26, n_100);
  and g219 (n_251, wc27, n_70);
  not gc27 (wc27, n_107);
  and g220 (n_252, wc28, n_227);
  not gc28 (wc28, n_246);
  and g221 (n_253, wc29, n_82);
  not gc29 (wc29, n_117);
  and g222 (n_148, wc30, n_228);
  not gc30 (wc30, n_247);
  and g223 (n_254, wc31, n_94);
  not gc31 (wc31, n_127);
  and g224 (n_255, wc32, n_129);
  not gc32 (wc32, n_148);
  or g225 (n_256, wc33, n_69);
  not gc33 (wc33, n_136);
  or g226 (n_257, n_229, wc34);
  not gc34 (wc34, n_136);
  or g227 (n_258, n_144, wc35);
  not gc35 (wc35, n_136);
  and g228 (n_259, wc36, n_88);
  not gc36 (wc36, n_149);
  and g229 (n_260, wc37, n_126);
  not gc37 (wc37, n_255);
  and g230 (n_261, n_254, wc38);
  not gc38 (wc38, n_157);
  or g231 (n_262, wc39, n_81);
  not gc39 (wc39, n_163);
  or g232 (n_263, n_230, wc40);
  not gc40 (wc40, n_163);
  or g233 (n_264, wc41, n_151);
  not gc41 (wc41, n_163);
endmodule

module add_unsigned_32_GENERIC(A, B, Z);
  input [15:0] A, B;
  output [15:0] Z;
  wire [15:0] A, B;
  wire [15:0] Z;
  add_unsigned_32_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_carry_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_unsigned_carry
  input [16:0] A, B;
  input CI;
  output [16:0] Z;
  wire [16:0] A, B;
  wire CI;
  wire [16:0] Z;
  wire n_53, n_54, n_55, n_56, n_57, n_59, n_61, n_62;
  wire n_63, n_64, n_66, n_67, n_68, n_69, n_70, n_72;
  wire n_73, n_74, n_75, n_76, n_78, n_79, n_80, n_81;
  wire n_82, n_84, n_85, n_86, n_87, n_88, n_90, n_91;
  wire n_92, n_93, n_94, n_96, n_97, n_98, n_99, n_100;
  wire n_102, n_103, n_106, n_108, n_109, n_110, n_112, n_114;
  wire n_119, n_120, n_122, n_124, n_129, n_130, n_132, n_134;
  wire n_139, n_142, n_147, n_151, n_152, n_154, n_158, n_160;
  wire n_162, n_164, n_166, n_169, n_176, n_178, n_181, n_182;
  wire n_184, n_185, n_187, n_188, n_189, n_191, n_196, n_200;
  wire n_202, n_205, n_209, n_211, n_214, n_217, n_220, n_222;
  wire n_225, n_228, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277;
  xor g1 (n_228, A[0], B[0]);
  nand g2 (n_53, A[0], B[0]);
  nand g3 (n_54, A[0], CI);
  nand g4 (n_55, B[0], CI);
  nand g5 (n_57, n_53, n_54, n_55);
  nor g6 (n_56, A[1], B[1]);
  nand g7 (n_59, A[1], B[1]);
  nor g8 (n_66, A[2], B[2]);
  nand g9 (n_61, A[2], B[2]);
  nor g10 (n_62, A[3], B[3]);
  nand g11 (n_63, A[3], B[3]);
  nor g12 (n_72, A[4], B[4]);
  nand g13 (n_67, A[4], B[4]);
  nor g14 (n_68, A[5], B[5]);
  nand g15 (n_69, A[5], B[5]);
  nor g16 (n_78, A[6], B[6]);
  nand g17 (n_73, A[6], B[6]);
  nor g18 (n_74, A[7], B[7]);
  nand g19 (n_75, A[7], B[7]);
  nor g20 (n_84, A[8], B[8]);
  nand g21 (n_79, A[8], B[8]);
  nor g22 (n_80, A[9], B[9]);
  nand g23 (n_81, A[9], B[9]);
  nor g24 (n_90, A[10], B[10]);
  nand g25 (n_85, A[10], B[10]);
  nor g26 (n_86, A[11], B[11]);
  nand g27 (n_87, A[11], B[11]);
  nor g28 (n_96, A[12], B[12]);
  nand g29 (n_91, A[12], B[12]);
  nor g30 (n_92, A[13], B[13]);
  nand g31 (n_93, A[13], B[13]);
  nor g32 (n_102, A[14], B[14]);
  nand g33 (n_97, A[14], B[14]);
  nor g34 (n_98, A[15], B[15]);
  nand g35 (n_99, A[15], B[15]);
  nor g36 (n_188, A[16], B[16]);
  nand g37 (n_191, A[16], B[16]);
  nand g40 (n_103, n_59, n_234);
  nor g41 (n_64, n_61, n_62);
  nor g44 (n_106, n_66, n_62);
  nor g45 (n_70, n_67, n_68);
  nor g48 (n_112, n_72, n_68);
  nor g49 (n_76, n_73, n_74);
  nor g52 (n_114, n_78, n_74);
  nor g53 (n_82, n_79, n_80);
  nor g56 (n_122, n_84, n_80);
  nor g57 (n_88, n_85, n_86);
  nor g60 (n_124, n_90, n_86);
  nor g61 (n_94, n_91, n_92);
  nor g64 (n_132, n_96, n_92);
  nor g65 (n_100, n_97, n_98);
  nor g68 (n_134, n_102, n_98);
  nand g71 (n_196, n_61, n_261);
  nand g72 (n_108, n_106, n_103);
  nand g73 (n_139, n_235, n_108);
  nor g74 (n_110, n_78, n_109);
  nand g83 (n_147, n_112, n_114);
  nor g84 (n_120, n_90, n_119);
  nand g93 (n_154, n_122, n_124);
  nor g94 (n_130, n_102, n_129);
  nand g103 (n_162, n_132, n_134);
  nand g106 (n_200, n_67, n_268);
  nand g107 (n_142, n_112, n_139);
  nand g108 (n_202, n_109, n_142);
  nand g111 (n_205, n_262, n_269);
  nand g114 (n_166, n_263, n_270);
  nor g115 (n_152, n_96, n_151);
  nor g118 (n_176, n_96, n_154);
  nor g124 (n_160, n_158, n_151);
  nor g127 (n_182, n_154, n_158);
  nor g128 (n_164, n_162, n_151);
  nor g131 (n_185, n_154, n_162);
  nand g134 (n_209, n_79, n_275);
  nand g135 (n_169, n_122, n_166);
  nand g136 (n_211, n_119, n_169);
  nand g139 (n_214, n_264, n_276);
  nand g142 (n_217, n_151, n_277);
  nand g143 (n_178, n_176, n_166);
  nand g144 (n_220, n_271, n_178);
  nand g145 (n_181, n_260, n_166);
  nand g146 (n_222, n_272, n_181);
  nand g147 (n_184, n_182, n_166);
  nand g148 (n_225, n_273, n_184);
  nand g149 (n_187, n_185, n_166);
  nand g150 (n_189, n_274, n_187);
  xnor g155 (Z[1], n_57, n_241);
  xnor g157 (Z[2], n_103, n_242);
  xnor g160 (Z[3], n_196, n_243);
  xnor g162 (Z[4], n_139, n_244);
  xnor g165 (Z[5], n_200, n_245);
  xnor g167 (Z[6], n_202, n_246);
  xnor g170 (Z[7], n_205, n_247);
  xnor g172 (Z[8], n_166, n_248);
  xnor g175 (Z[9], n_209, n_249);
  xnor g177 (Z[10], n_211, n_250);
  xnor g180 (Z[11], n_214, n_251);
  xnor g183 (Z[12], n_217, n_252);
  xnor g186 (Z[13], n_220, n_253);
  xnor g188 (Z[14], n_222, n_254);
  xnor g191 (Z[15], n_225, n_255);
  xnor g193 (Z[16], n_189, n_256);
  xor g194 (Z[0], CI, n_228);
  or g195 (n_234, n_56, wc);
  not gc (wc, n_57);
  and g196 (n_235, wc0, n_63);
  not gc0 (wc0, n_64);
  and g197 (n_109, wc1, n_69);
  not gc1 (wc1, n_70);
  and g198 (n_236, wc2, n_75);
  not gc2 (wc2, n_76);
  and g199 (n_119, wc3, n_81);
  not gc3 (wc3, n_82);
  and g200 (n_237, wc4, n_87);
  not gc4 (wc4, n_88);
  and g201 (n_129, wc5, n_93);
  not gc5 (wc5, n_94);
  and g202 (n_238, wc6, n_99);
  not gc6 (wc6, n_100);
  or g203 (n_239, wc7, n_78);
  not gc7 (wc7, n_112);
  or g204 (n_240, wc8, n_90);
  not gc8 (wc8, n_122);
  or g205 (n_158, wc9, n_102);
  not gc9 (wc9, n_132);
  or g206 (n_241, wc10, n_56);
  not gc10 (wc10, n_59);
  or g207 (n_242, wc11, n_66);
  not gc11 (wc11, n_61);
  or g208 (n_243, wc12, n_62);
  not gc12 (wc12, n_63);
  or g209 (n_244, wc13, n_72);
  not gc13 (wc13, n_67);
  or g210 (n_245, wc14, n_68);
  not gc14 (wc14, n_69);
  or g211 (n_246, wc15, n_78);
  not gc15 (wc15, n_73);
  or g212 (n_247, wc16, n_74);
  not gc16 (wc16, n_75);
  or g213 (n_248, wc17, n_84);
  not gc17 (wc17, n_79);
  or g214 (n_249, wc18, n_80);
  not gc18 (wc18, n_81);
  or g215 (n_250, wc19, n_90);
  not gc19 (wc19, n_85);
  or g216 (n_251, wc20, n_86);
  not gc20 (wc20, n_87);
  or g217 (n_252, wc21, n_96);
  not gc21 (wc21, n_91);
  or g218 (n_253, wc22, n_92);
  not gc22 (wc22, n_93);
  or g219 (n_254, wc23, n_102);
  not gc23 (wc23, n_97);
  or g220 (n_255, wc24, n_98);
  not gc24 (wc24, n_99);
  or g221 (n_256, wc25, n_188);
  not gc25 (wc25, n_191);
  and g222 (n_257, wc26, n_114);
  not gc26 (wc26, n_109);
  and g223 (n_258, wc27, n_124);
  not gc27 (wc27, n_119);
  and g224 (n_259, wc28, n_134);
  not gc28 (wc28, n_129);
  and g225 (n_260, wc29, n_132);
  not gc29 (wc29, n_154);
  or g226 (n_261, wc30, n_66);
  not gc30 (wc30, n_103);
  and g227 (n_262, wc31, n_73);
  not gc31 (wc31, n_110);
  and g228 (n_263, wc32, n_236);
  not gc32 (wc32, n_257);
  and g229 (n_264, wc33, n_85);
  not gc33 (wc33, n_120);
  and g230 (n_151, wc34, n_237);
  not gc34 (wc34, n_258);
  and g231 (n_265, wc35, n_97);
  not gc35 (wc35, n_130);
  and g232 (n_266, wc36, n_238);
  not gc36 (wc36, n_259);
  and g233 (n_267, wc37, n_132);
  not gc37 (wc37, n_151);
  or g234 (n_268, wc38, n_72);
  not gc38 (wc38, n_139);
  or g235 (n_269, n_239, wc39);
  not gc39 (wc39, n_139);
  or g236 (n_270, n_147, wc40);
  not gc40 (wc40, n_139);
  and g237 (n_271, wc41, n_91);
  not gc41 (wc41, n_152);
  and g238 (n_272, wc42, n_129);
  not gc42 (wc42, n_267);
  and g239 (n_273, n_265, wc43);
  not gc43 (wc43, n_160);
  and g240 (n_274, n_266, wc44);
  not gc44 (wc44, n_164);
  or g241 (n_275, wc45, n_84);
  not gc45 (wc45, n_166);
  or g242 (n_276, n_240, wc46);
  not gc46 (wc46, n_166);
  or g243 (n_277, wc47, n_154);
  not gc47 (wc47, n_166);
endmodule

module add_unsigned_carry_GENERIC(A, B, CI, Z);
  input [16:0] A, B;
  input CI;
  output [16:0] Z;
  wire [16:0] A, B;
  wire CI;
  wire [16:0] Z;
  add_unsigned_carry_GENERIC_REAL g1(.A (A), .B (B), .CI (CI), .Z (Z));
endmodule

module bmux_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [16:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  or g18 (z[16], wc, wc1);
  and gc1 (wc1, in_1[16], ctl);
  and gc0 (wc, in_0[16], wc0);
  not gc (wc0, ctl);
  or g19 (z[15], wc2, wc4);
  and gc4 (wc4, in_1[15], ctl);
  and gc3 (wc2, in_0[15], wc3);
  not gc2 (wc3, ctl);
  or g20 (z[14], wc5, wc7);
  and gc7 (wc7, in_1[14], ctl);
  and gc6 (wc5, in_0[14], wc6);
  not gc5 (wc6, ctl);
  or g21 (z[13], wc8, wc10);
  and gc10 (wc10, in_1[13], ctl);
  and gc9 (wc8, in_0[13], wc9);
  not gc8 (wc9, ctl);
  or g22 (z[12], wc11, wc13);
  and gc13 (wc13, in_1[12], ctl);
  and gc12 (wc11, in_0[12], wc12);
  not gc11 (wc12, ctl);
  or g23 (z[11], wc14, wc16);
  and gc16 (wc16, in_1[11], ctl);
  and gc15 (wc14, in_0[11], wc15);
  not gc14 (wc15, ctl);
  or g24 (z[10], wc17, wc19);
  and gc19 (wc19, in_1[10], ctl);
  and gc18 (wc17, in_0[10], wc18);
  not gc17 (wc18, ctl);
  or g25 (z[9], wc20, wc22);
  and gc22 (wc22, in_1[9], ctl);
  and gc21 (wc20, in_0[9], wc21);
  not gc20 (wc21, ctl);
  or g26 (z[8], wc23, wc25);
  and gc25 (wc25, in_1[8], ctl);
  and gc24 (wc23, in_0[8], wc24);
  not gc23 (wc24, ctl);
  or g27 (z[7], wc26, wc28);
  and gc28 (wc28, in_1[7], ctl);
  and gc27 (wc26, in_0[7], wc27);
  not gc26 (wc27, ctl);
  or g28 (z[6], wc29, wc31);
  and gc31 (wc31, in_1[6], ctl);
  and gc30 (wc29, in_0[6], wc30);
  not gc29 (wc30, ctl);
  or g29 (z[5], wc32, wc34);
  and gc34 (wc34, in_1[5], ctl);
  and gc33 (wc32, in_0[5], wc33);
  not gc32 (wc33, ctl);
  or g30 (z[4], wc35, wc37);
  and gc37 (wc37, in_1[4], ctl);
  and gc36 (wc35, in_0[4], wc36);
  not gc35 (wc36, ctl);
  or g31 (z[3], wc38, wc40);
  and gc40 (wc40, in_1[3], ctl);
  and gc39 (wc38, in_0[3], wc39);
  not gc38 (wc39, ctl);
  or g32 (z[2], wc41, wc43);
  and gc43 (wc43, in_1[2], ctl);
  and gc42 (wc41, in_0[2], wc42);
  not gc41 (wc42, ctl);
  or g33 (z[1], wc44, wc46);
  and gc46 (wc46, in_1[1], ctl);
  and gc45 (wc44, in_0[1], wc45);
  not gc44 (wc45, ctl);
  or g34 (z[0], wc47, wc49);
  and gc49 (wc49, in_1[0], ctl);
  and gc48 (wc47, in_0[0], wc48);
  not gc47 (wc48, ctl);
endmodule

module bmux_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  bmux_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1), .z (z));
endmodule

module bmux_1_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [16:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  or g18 (z[16], wc, wc1);
  and gc1 (wc1, in_1[16], ctl);
  and gc0 (wc, in_0[16], wc0);
  not gc (wc0, ctl);
  or g19 (z[15], wc2, wc4);
  and gc4 (wc4, in_1[15], ctl);
  and gc3 (wc2, in_0[15], wc3);
  not gc2 (wc3, ctl);
  or g20 (z[14], wc5, wc7);
  and gc7 (wc7, in_1[14], ctl);
  and gc6 (wc5, in_0[14], wc6);
  not gc5 (wc6, ctl);
  or g21 (z[13], wc8, wc10);
  and gc10 (wc10, in_1[13], ctl);
  and gc9 (wc8, in_0[13], wc9);
  not gc8 (wc9, ctl);
  or g22 (z[12], wc11, wc13);
  and gc13 (wc13, in_1[12], ctl);
  and gc12 (wc11, in_0[12], wc12);
  not gc11 (wc12, ctl);
  or g23 (z[11], wc14, wc16);
  and gc16 (wc16, in_1[11], ctl);
  and gc15 (wc14, in_0[11], wc15);
  not gc14 (wc15, ctl);
  or g24 (z[10], wc17, wc19);
  and gc19 (wc19, in_1[10], ctl);
  and gc18 (wc17, in_0[10], wc18);
  not gc17 (wc18, ctl);
  or g25 (z[9], wc20, wc22);
  and gc22 (wc22, in_1[9], ctl);
  and gc21 (wc20, in_0[9], wc21);
  not gc20 (wc21, ctl);
  or g26 (z[8], wc23, wc25);
  and gc25 (wc25, in_1[8], ctl);
  and gc24 (wc23, in_0[8], wc24);
  not gc23 (wc24, ctl);
  or g27 (z[7], wc26, wc28);
  and gc28 (wc28, in_1[7], ctl);
  and gc27 (wc26, in_0[7], wc27);
  not gc26 (wc27, ctl);
  or g28 (z[6], wc29, wc31);
  and gc31 (wc31, in_1[6], ctl);
  and gc30 (wc29, in_0[6], wc30);
  not gc29 (wc30, ctl);
  or g29 (z[5], wc32, wc34);
  and gc34 (wc34, in_1[5], ctl);
  and gc33 (wc32, in_0[5], wc33);
  not gc32 (wc33, ctl);
  or g30 (z[4], wc35, wc37);
  and gc37 (wc37, in_1[4], ctl);
  and gc36 (wc35, in_0[4], wc36);
  not gc35 (wc36, ctl);
  or g31 (z[3], wc38, wc40);
  and gc40 (wc40, in_1[3], ctl);
  and gc39 (wc38, in_0[3], wc39);
  not gc38 (wc39, ctl);
  or g32 (z[2], wc41, wc43);
  and gc43 (wc43, in_1[2], ctl);
  and gc42 (wc41, in_0[2], wc42);
  not gc41 (wc42, ctl);
  or g33 (z[1], wc44, wc46);
  and gc46 (wc46, in_1[1], ctl);
  and gc45 (wc44, in_0[1], wc45);
  not gc44 (wc45, ctl);
  or g34 (z[0], wc47, wc49);
  and gc49 (wc49, in_1[0], ctl);
  and gc48 (wc47, in_0[0], wc48);
  not gc47 (wc48, ctl);
endmodule

module bmux_1_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  bmux_1_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1), .z
       (z));
endmodule

module csa_tree_GENERIC_REAL(in_0, in_1, out_0, out_1);
// synthesis_equation "assign out_0 = ( in_0 * in_1 )  ; assign out_1 = 16'b0;"
  input [7:0] in_0, in_1;
  output [15:0] out_0, out_1;
  wire [7:0] in_0, in_1;
  wire [15:0] out_0, out_1;
  wire n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305;
  assign out_1[0] = 1'b0;
  assign out_1[15] = 1'b0;
  assign out_0[15] = 1'b0;
  and g1 (out_0[0], in_0[0], in_1[0]);
  and g2 (out_0[1], in_0[1], in_1[0]);
  and g3 (n_17, in_0[2], in_1[0]);
  and g4 (n_19, in_0[3], in_1[0]);
  and g5 (n_24, in_0[4], in_1[0]);
  and g6 (n_32, in_0[5], in_1[0]);
  and g7 (n_43, in_0[6], in_1[0]);
  and g8 (n_57, in_0[7], in_1[0]);
  and g9 (out_1[1], in_0[0], in_1[1]);
  and g10 (out_0[2], in_0[1], in_1[1]);
  and g11 (n_20, in_0[2], in_1[1]);
  and g12 (n_25, in_0[3], in_1[1]);
  and g13 (n_33, in_0[4], in_1[1]);
  and g14 (n_44, in_0[5], in_1[1]);
  and g15 (n_58, in_0[6], in_1[1]);
  and g16 (n_74, in_0[7], in_1[1]);
  and g17 (n_18, in_0[0], in_1[2]);
  and g18 (n_22, in_0[1], in_1[2]);
  and g19 (n_28, in_0[2], in_1[2]);
  and g20 (n_36, in_0[3], in_1[2]);
  and g21 (n_47, in_0[4], in_1[2]);
  and g22 (n_62, in_0[5], in_1[2]);
  and g23 (n_75, in_0[6], in_1[2]);
  and g24 (n_91, in_0[7], in_1[2]);
  and g25 (n_21, in_0[0], in_1[3]);
  and g26 (n_26, in_0[1], in_1[3]);
  and g27 (n_34, in_0[2], in_1[3]);
  and g28 (n_45, in_0[3], in_1[3]);
  and g29 (n_59, in_0[4], in_1[3]);
  and g30 (n_78, in_0[5], in_1[3]);
  and g31 (n_92, in_0[6], in_1[3]);
  and g32 (n_106, in_0[7], in_1[3]);
  and g33 (n_27, in_0[0], in_1[4]);
  and g34 (n_35, in_0[1], in_1[4]);
  and g35 (n_46, in_0[2], in_1[4]);
  and g36 (n_61, in_0[3], in_1[4]);
  and g37 (n_76, in_0[4], in_1[4]);
  and g38 (n_95, in_0[5], in_1[4]);
  and g39 (n_107, in_0[6], in_1[4]);
  and g40 (n_118, in_0[7], in_1[4]);
  and g41 (n_37, in_0[0], in_1[5]);
  and g42 (n_48, in_0[1], in_1[5]);
  and g43 (n_63, in_0[2], in_1[5]);
  and g44 (n_77, in_0[3], in_1[5]);
  and g45 (n_93, in_0[4], in_1[5]);
  and g46 (n_110, in_0[5], in_1[5]);
  and g47 (n_119, in_0[6], in_1[5]);
  and g48 (n_127, in_0[7], in_1[5]);
  and g49 (n_49, in_0[0], in_1[6]);
  and g50 (n_64, in_0[1], in_1[6]);
  and g51 (n_79, in_0[2], in_1[6]);
  and g52 (n_94, in_0[3], in_1[6]);
  and g53 (n_108, in_0[4], in_1[6]);
  and g54 (n_121, in_0[5], in_1[6]);
  and g55 (n_128, in_0[6], in_1[6]);
  and g56 (n_133, in_0[7], in_1[6]);
  and g57 (n_60, in_0[0], in_1[7]);
  and g58 (n_80, in_0[1], in_1[7]);
  and g59 (n_96, in_0[2], in_1[7]);
  and g60 (n_109, in_0[3], in_1[7]);
  and g61 (n_120, in_0[4], in_1[7]);
  and g62 (n_129, in_0[5], in_1[7]);
  and g63 (n_134, in_0[6], in_1[7]);
  and g64 (out_0[14], in_0[7], in_1[7]);
  xor g107 (out_1[2], n_17, n_18);
  and g108 (out_0[3], n_17, n_18);
  xor g109 (n_23, n_19, n_20);
  and g110 (n_30, n_19, n_20);
  xor g111 (n_166, n_21, n_22);
  xor g112 (out_1[3], n_166, n_23);
  nand g113 (n_167, n_21, n_22);
  nand g114 (n_168, n_23, n_22);
  nand g115 (n_169, n_21, n_23);
  nand g116 (out_0[4], n_167, n_168, n_169);
  xor g117 (n_29, n_24, n_25);
  and g118 (n_39, n_24, n_25);
  xor g119 (n_170, n_26, n_27);
  xor g120 (n_31, n_170, n_28);
  nand g121 (n_171, n_26, n_27);
  nand g122 (n_172, n_28, n_27);
  nand g123 (n_173, n_26, n_28);
  nand g124 (n_40, n_171, n_172, n_173);
  xor g125 (n_174, n_29, n_30);
  xor g126 (out_1[4], n_174, n_31);
  nand g127 (n_175, n_29, n_30);
  nand g128 (n_176, n_31, n_30);
  nand g129 (n_177, n_29, n_31);
  nand g130 (out_0[5], n_175, n_176, n_177);
  xor g131 (n_38, n_32, n_33);
  and g132 (n_50, n_32, n_33);
  xor g133 (n_178, n_34, n_35);
  xor g134 (n_41, n_178, n_36);
  nand g135 (n_179, n_34, n_35);
  nand g136 (n_180, n_36, n_35);
  nand g137 (n_181, n_34, n_36);
  nand g138 (n_52, n_179, n_180, n_181);
  xor g139 (n_182, n_37, n_38);
  xor g140 (n_42, n_182, n_39);
  nand g141 (n_183, n_37, n_38);
  nand g142 (n_184, n_39, n_38);
  nand g143 (n_185, n_37, n_39);
  nand g144 (n_54, n_183, n_184, n_185);
  xor g145 (n_186, n_40, n_41);
  xor g146 (out_1[5], n_186, n_42);
  nand g147 (n_187, n_40, n_41);
  nand g148 (n_188, n_42, n_41);
  nand g149 (n_189, n_40, n_42);
  nand g150 (out_0[6], n_187, n_188, n_189);
  xor g151 (n_51, n_43, n_44);
  and g152 (n_65, n_43, n_44);
  xor g153 (n_190, n_45, n_46);
  xor g154 (n_53, n_190, n_47);
  nand g155 (n_191, n_45, n_46);
  nand g156 (n_192, n_47, n_46);
  nand g157 (n_193, n_45, n_47);
  nand g158 (n_67, n_191, n_192, n_193);
  xor g159 (n_194, n_48, n_49);
  xor g160 (n_55, n_194, n_50);
  nand g161 (n_195, n_48, n_49);
  nand g162 (n_196, n_50, n_49);
  nand g163 (n_197, n_48, n_50);
  nand g164 (n_70, n_195, n_196, n_197);
  xor g165 (n_198, n_51, n_52);
  xor g166 (n_56, n_198, n_53);
  nand g167 (n_199, n_51, n_52);
  nand g168 (n_200, n_53, n_52);
  nand g169 (n_201, n_51, n_53);
  nand g170 (n_72, n_199, n_200, n_201);
  xor g171 (n_202, n_54, n_55);
  xor g172 (out_1[6], n_202, n_56);
  nand g173 (n_203, n_54, n_55);
  nand g174 (n_204, n_56, n_55);
  nand g175 (n_205, n_54, n_56);
  nand g176 (out_0[7], n_203, n_204, n_205);
  xor g177 (n_66, n_57, n_58);
  and g178 (n_82, n_57, n_58);
  xor g179 (n_206, n_59, n_60);
  xor g180 (n_69, n_206, n_61);
  nand g181 (n_207, n_59, n_60);
  nand g182 (n_208, n_61, n_60);
  nand g183 (n_209, n_59, n_61);
  nand g184 (n_83, n_207, n_208, n_209);
  xor g185 (n_210, n_62, n_63);
  xor g186 (n_68, n_210, n_64);
  nand g187 (n_211, n_62, n_63);
  nand g188 (n_212, n_64, n_63);
  nand g189 (n_213, n_62, n_64);
  nand g190 (n_84, n_211, n_212, n_213);
  xor g191 (n_214, n_65, n_66);
  xor g192 (n_71, n_214, n_67);
  nand g193 (n_215, n_65, n_66);
  nand g194 (n_216, n_67, n_66);
  nand g195 (n_217, n_65, n_67);
  nand g196 (n_87, n_215, n_216, n_217);
  xor g197 (n_218, n_68, n_69);
  xor g198 (n_73, n_218, n_70);
  nand g199 (n_219, n_68, n_69);
  nand g200 (n_220, n_70, n_69);
  nand g201 (n_221, n_68, n_70);
  nand g202 (n_89, n_219, n_220, n_221);
  xor g203 (n_222, n_71, n_72);
  xor g204 (out_1[7], n_222, n_73);
  nand g205 (n_223, n_71, n_72);
  nand g206 (n_224, n_73, n_72);
  nand g207 (n_225, n_71, n_73);
  nand g208 (out_0[8], n_223, n_224, n_225);
  xor g209 (n_81, n_74, n_75);
  and g210 (n_97, n_74, n_75);
  xor g211 (n_226, n_76, n_77);
  xor g212 (n_85, n_226, n_78);
  nand g213 (n_227, n_76, n_77);
  nand g214 (n_228, n_78, n_77);
  nand g215 (n_229, n_76, n_78);
  nand g216 (n_98, n_227, n_228, n_229);
  xor g217 (n_230, n_79, n_80);
  xor g218 (n_86, n_230, n_81);
  nand g219 (n_231, n_79, n_80);
  nand g220 (n_232, n_81, n_80);
  nand g221 (n_233, n_79, n_81);
  nand g222 (n_101, n_231, n_232, n_233);
  xor g223 (n_234, n_82, n_83);
  xor g224 (n_88, n_234, n_84);
  nand g225 (n_235, n_82, n_83);
  nand g226 (n_236, n_84, n_83);
  nand g227 (n_237, n_82, n_84);
  nand g228 (n_102, n_235, n_236, n_237);
  xor g229 (n_238, n_85, n_86);
  xor g230 (n_90, n_238, n_87);
  nand g231 (n_239, n_85, n_86);
  nand g232 (n_240, n_87, n_86);
  nand g233 (n_241, n_85, n_87);
  nand g234 (n_105, n_239, n_240, n_241);
  xor g235 (n_242, n_88, n_89);
  xor g236 (out_1[8], n_242, n_90);
  nand g237 (n_243, n_88, n_89);
  nand g238 (n_244, n_90, n_89);
  nand g239 (n_245, n_88, n_90);
  nand g240 (out_0[9], n_243, n_244, n_245);
  xor g241 (n_246, n_91, n_92);
  xor g242 (n_100, n_246, n_93);
  nand g243 (n_247, n_91, n_92);
  nand g244 (n_248, n_93, n_92);
  nand g245 (n_249, n_91, n_93);
  nand g246 (n_112, n_247, n_248, n_249);
  xor g247 (n_250, n_94, n_95);
  xor g248 (n_99, n_250, n_96);
  nand g249 (n_251, n_94, n_95);
  nand g250 (n_252, n_96, n_95);
  nand g251 (n_253, n_94, n_96);
  nand g252 (n_111, n_251, n_252, n_253);
  xor g253 (n_254, n_97, n_98);
  xor g254 (n_103, n_254, n_99);
  nand g255 (n_255, n_97, n_98);
  nand g256 (n_256, n_99, n_98);
  nand g257 (n_257, n_97, n_99);
  nand g258 (n_115, n_255, n_256, n_257);
  xor g259 (n_258, n_100, n_101);
  xor g260 (n_104, n_258, n_102);
  nand g261 (n_259, n_100, n_101);
  nand g262 (n_260, n_102, n_101);
  nand g263 (n_261, n_100, n_102);
  nand g264 (n_117, n_259, n_260, n_261);
  xor g265 (n_262, n_103, n_104);
  xor g266 (out_1[9], n_262, n_105);
  nand g267 (n_263, n_103, n_104);
  nand g268 (n_264, n_105, n_104);
  nand g269 (n_265, n_103, n_105);
  nand g270 (out_0[10], n_263, n_264, n_265);
  xor g271 (n_266, n_106, n_107);
  xor g272 (n_113, n_266, n_108);
  nand g273 (n_267, n_106, n_107);
  nand g274 (n_268, n_108, n_107);
  nand g275 (n_269, n_106, n_108);
  nand g276 (n_122, n_267, n_268, n_269);
  xor g277 (n_270, n_109, n_110);
  xor g278 (n_114, n_270, n_111);
  nand g279 (n_271, n_109, n_110);
  nand g280 (n_272, n_111, n_110);
  nand g281 (n_273, n_109, n_111);
  nand g282 (n_124, n_271, n_272, n_273);
  xor g283 (n_274, n_112, n_113);
  xor g284 (n_116, n_274, n_114);
  nand g285 (n_275, n_112, n_113);
  nand g286 (n_276, n_114, n_113);
  nand g287 (n_277, n_112, n_114);
  nand g288 (n_126, n_275, n_276, n_277);
  xor g289 (n_278, n_115, n_116);
  xor g290 (out_1[10], n_278, n_117);
  nand g291 (n_279, n_115, n_116);
  nand g292 (n_280, n_117, n_116);
  nand g293 (n_281, n_115, n_117);
  nand g294 (out_0[11], n_279, n_280, n_281);
  xor g295 (n_282, n_118, n_119);
  xor g296 (n_123, n_282, n_120);
  nand g297 (n_283, n_118, n_119);
  nand g298 (n_284, n_120, n_119);
  nand g299 (n_285, n_118, n_120);
  nand g300 (n_130, n_283, n_284, n_285);
  xor g301 (n_286, n_121, n_122);
  xor g302 (n_125, n_286, n_123);
  nand g303 (n_287, n_121, n_122);
  nand g304 (n_288, n_123, n_122);
  nand g305 (n_289, n_121, n_123);
  nand g306 (n_132, n_287, n_288, n_289);
  xor g307 (n_290, n_124, n_125);
  xor g308 (out_1[11], n_290, n_126);
  nand g309 (n_291, n_124, n_125);
  nand g310 (n_292, n_126, n_125);
  nand g311 (n_293, n_124, n_126);
  nand g312 (out_1[12], n_291, n_292, n_293);
  xor g313 (n_294, n_127, n_128);
  xor g314 (n_131, n_294, n_129);
  nand g315 (n_295, n_127, n_128);
  nand g316 (n_296, n_129, n_128);
  nand g317 (n_297, n_127, n_129);
  nand g318 (n_135, n_295, n_296, n_297);
  xor g319 (n_298, n_130, n_131);
  xor g320 (out_0[12], n_298, n_132);
  nand g321 (n_299, n_130, n_131);
  nand g322 (n_300, n_132, n_131);
  nand g323 (n_301, n_130, n_132);
  nand g324 (out_1[13], n_299, n_300, n_301);
  xor g325 (n_302, n_133, n_134);
  xor g326 (out_0[13], n_302, n_135);
  nand g327 (n_303, n_133, n_134);
  nand g328 (n_304, n_135, n_134);
  nand g329 (n_305, n_133, n_135);
  nand g330 (out_1[14], n_303, n_304, n_305);
endmodule

module csa_tree_GENERIC(in_0, in_1, out_0, out_1);
  input [7:0] in_0, in_1;
  output [15:0] out_0, out_1;
  wire [7:0] in_0, in_1;
  wire [15:0] out_0, out_1;
  csa_tree_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .out_0 (out_0),
       .out_1 (out_1));
endmodule

module csa_tree_112_GENERIC_REAL(in_0, in_1, in_2, in_3, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( in_0 + in_1 ) + ( in_2 + in_3 ) )  ; assign out_1 = 17'b0;"
  input [15:0] in_0, in_1, in_2, in_3;
  output [16:0] out_0, out_1;
  wire [15:0] in_0, in_1, in_2, in_3;
  wire [16:0] out_0, out_1;
  wire n_8, n_13, n_14, n_19, n_20, n_25, n_26, n_31;
  wire n_32, n_37, n_38, n_43, n_44, n_49, n_50, n_55;
  wire n_56, n_61, n_62, n_67, n_68, n_73, n_74, n_79;
  wire n_80, n_85, n_86, n_91, n_92, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246;
  assign out_0[0] = in_1[0];
  xor g1 (n_127, in_0[0], in_3[0]);
  xor g32 (out_1[0], n_127, in_2[0]);
  nand g33 (n_128, in_0[0], in_3[0]);
  nand g34 (n_129, in_2[0], in_3[0]);
  nand g35 (n_130, in_0[0], in_2[0]);
  nand g36 (out_0[1], n_128, n_129, n_130);
  xor g37 (n_8, in_0[1], in_1[1]);
  and g2 (n_13, in_0[1], in_1[1]);
  xor g38 (n_131, in_3[1], in_2[1]);
  xor g39 (out_1[1], n_131, n_8);
  nand g3 (n_132, in_3[1], in_2[1]);
  nand g40 (n_133, n_8, in_2[1]);
  nand g41 (n_134, in_3[1], n_8);
  nand g42 (out_0[2], n_132, n_133, n_134);
  xor g43 (n_135, in_0[2], in_1[2]);
  xor g44 (n_14, n_135, in_3[2]);
  nand g45 (n_136, in_0[2], in_1[2]);
  nand g4 (n_137, in_3[2], in_1[2]);
  nand g46 (n_138, in_0[2], in_3[2]);
  nand g47 (n_19, n_136, n_137, n_138);
  xor g48 (n_139, in_2[2], n_13);
  xor g49 (out_1[2], n_139, n_14);
  nand g50 (n_140, in_2[2], n_13);
  nand g51 (n_141, n_14, n_13);
  nand g5 (n_142, in_2[2], n_14);
  nand g52 (out_0[3], n_140, n_141, n_142);
  xor g53 (n_143, in_0[3], in_1[3]);
  xor g54 (n_20, n_143, in_3[3]);
  nand g55 (n_144, in_0[3], in_1[3]);
  nand g56 (n_145, in_3[3], in_1[3]);
  nand g57 (n_146, in_0[3], in_3[3]);
  nand g6 (n_25, n_144, n_145, n_146);
  xor g58 (n_147, in_2[3], n_19);
  xor g59 (out_1[3], n_147, n_20);
  nand g60 (n_148, in_2[3], n_19);
  nand g61 (n_149, n_20, n_19);
  nand g62 (n_150, in_2[3], n_20);
  nand g63 (out_0[4], n_148, n_149, n_150);
  xor g64 (n_151, in_0[4], in_1[4]);
  xor g65 (n_26, n_151, in_3[4]);
  nand g66 (n_152, in_0[4], in_1[4]);
  nand g67 (n_153, in_3[4], in_1[4]);
  nand g68 (n_154, in_0[4], in_3[4]);
  nand g69 (n_31, n_152, n_153, n_154);
  xor g70 (n_155, in_2[4], n_25);
  xor g71 (out_1[4], n_155, n_26);
  nand g72 (n_156, in_2[4], n_25);
  nand g73 (n_157, n_26, n_25);
  nand g74 (n_158, in_2[4], n_26);
  nand g75 (out_0[5], n_156, n_157, n_158);
  xor g76 (n_159, in_0[5], in_1[5]);
  xor g77 (n_32, n_159, in_3[5]);
  nand g78 (n_160, in_0[5], in_1[5]);
  nand g79 (n_161, in_3[5], in_1[5]);
  nand g80 (n_162, in_0[5], in_3[5]);
  nand g81 (n_37, n_160, n_161, n_162);
  xor g82 (n_163, in_2[5], n_31);
  xor g83 (out_1[5], n_163, n_32);
  nand g84 (n_164, in_2[5], n_31);
  nand g85 (n_165, n_32, n_31);
  nand g86 (n_166, in_2[5], n_32);
  nand g87 (out_0[6], n_164, n_165, n_166);
  xor g88 (n_167, in_0[6], in_1[6]);
  xor g89 (n_38, n_167, in_3[6]);
  nand g90 (n_168, in_0[6], in_1[6]);
  nand g91 (n_169, in_3[6], in_1[6]);
  nand g92 (n_170, in_0[6], in_3[6]);
  nand g93 (n_43, n_168, n_169, n_170);
  xor g94 (n_171, in_2[6], n_37);
  xor g95 (out_1[6], n_171, n_38);
  nand g96 (n_172, in_2[6], n_37);
  nand g97 (n_173, n_38, n_37);
  nand g98 (n_174, in_2[6], n_38);
  nand g99 (out_0[7], n_172, n_173, n_174);
  xor g100 (n_175, in_0[7], in_1[7]);
  xor g101 (n_44, n_175, in_3[7]);
  nand g102 (n_176, in_0[7], in_1[7]);
  nand g103 (n_177, in_3[7], in_1[7]);
  nand g104 (n_178, in_0[7], in_3[7]);
  nand g105 (n_49, n_176, n_177, n_178);
  xor g106 (n_179, in_2[7], n_43);
  xor g107 (out_1[7], n_179, n_44);
  nand g108 (n_180, in_2[7], n_43);
  nand g109 (n_181, n_44, n_43);
  nand g110 (n_182, in_2[7], n_44);
  nand g111 (out_0[8], n_180, n_181, n_182);
  xor g112 (n_183, in_0[8], in_1[8]);
  xor g113 (n_50, n_183, in_3[8]);
  nand g114 (n_184, in_0[8], in_1[8]);
  nand g115 (n_185, in_3[8], in_1[8]);
  nand g116 (n_186, in_0[8], in_3[8]);
  nand g117 (n_55, n_184, n_185, n_186);
  xor g118 (n_187, in_2[8], n_49);
  xor g119 (out_1[8], n_187, n_50);
  nand g120 (n_188, in_2[8], n_49);
  nand g121 (n_189, n_50, n_49);
  nand g122 (n_190, in_2[8], n_50);
  nand g123 (out_0[9], n_188, n_189, n_190);
  xor g124 (n_191, in_0[9], in_1[9]);
  xor g125 (n_56, n_191, in_3[9]);
  nand g126 (n_192, in_0[9], in_1[9]);
  nand g127 (n_193, in_3[9], in_1[9]);
  nand g128 (n_194, in_0[9], in_3[9]);
  nand g129 (n_61, n_192, n_193, n_194);
  xor g130 (n_195, in_2[9], n_55);
  xor g131 (out_1[9], n_195, n_56);
  nand g132 (n_196, in_2[9], n_55);
  nand g133 (n_197, n_56, n_55);
  nand g134 (n_198, in_2[9], n_56);
  nand g135 (out_0[10], n_196, n_197, n_198);
  xor g136 (n_199, in_0[10], in_1[10]);
  xor g137 (n_62, n_199, in_3[10]);
  nand g138 (n_200, in_0[10], in_1[10]);
  nand g139 (n_201, in_3[10], in_1[10]);
  nand g140 (n_202, in_0[10], in_3[10]);
  nand g141 (n_67, n_200, n_201, n_202);
  xor g142 (n_203, in_2[10], n_61);
  xor g143 (out_1[10], n_203, n_62);
  nand g144 (n_204, in_2[10], n_61);
  nand g145 (n_205, n_62, n_61);
  nand g146 (n_206, in_2[10], n_62);
  nand g147 (out_0[11], n_204, n_205, n_206);
  xor g148 (n_207, in_0[11], in_1[11]);
  xor g149 (n_68, n_207, in_3[11]);
  nand g150 (n_208, in_0[11], in_1[11]);
  nand g151 (n_209, in_3[11], in_1[11]);
  nand g152 (n_210, in_0[11], in_3[11]);
  nand g153 (n_73, n_208, n_209, n_210);
  xor g154 (n_211, in_2[11], n_67);
  xor g155 (out_1[11], n_211, n_68);
  nand g156 (n_212, in_2[11], n_67);
  nand g157 (n_213, n_68, n_67);
  nand g158 (n_214, in_2[11], n_68);
  nand g159 (out_0[12], n_212, n_213, n_214);
  xor g160 (n_215, in_0[12], in_1[12]);
  xor g161 (n_74, n_215, in_3[12]);
  nand g162 (n_216, in_0[12], in_1[12]);
  nand g163 (n_217, in_3[12], in_1[12]);
  nand g164 (n_218, in_0[12], in_3[12]);
  nand g165 (n_79, n_216, n_217, n_218);
  xor g166 (n_219, in_2[12], n_73);
  xor g167 (out_1[12], n_219, n_74);
  nand g168 (n_220, in_2[12], n_73);
  nand g169 (n_221, n_74, n_73);
  nand g170 (n_222, in_2[12], n_74);
  nand g171 (out_0[13], n_220, n_221, n_222);
  xor g172 (n_223, in_0[13], in_1[13]);
  xor g173 (n_80, n_223, in_3[13]);
  nand g174 (n_224, in_0[13], in_1[13]);
  nand g175 (n_225, in_3[13], in_1[13]);
  nand g176 (n_226, in_0[13], in_3[13]);
  nand g177 (n_85, n_224, n_225, n_226);
  xor g178 (n_227, in_2[13], n_79);
  xor g179 (out_1[13], n_227, n_80);
  nand g180 (n_228, in_2[13], n_79);
  nand g181 (n_229, n_80, n_79);
  nand g182 (n_230, in_2[13], n_80);
  nand g183 (out_0[14], n_228, n_229, n_230);
  xor g184 (n_231, in_0[14], in_1[14]);
  xor g185 (n_86, n_231, in_3[14]);
  nand g186 (n_232, in_0[14], in_1[14]);
  nand g187 (n_233, in_3[14], in_1[14]);
  nand g188 (n_234, in_0[14], in_3[14]);
  nand g189 (n_91, n_232, n_233, n_234);
  xor g190 (n_235, in_2[14], n_85);
  xor g191 (out_1[14], n_235, n_86);
  nand g192 (n_236, in_2[14], n_85);
  nand g193 (n_237, n_86, n_85);
  nand g194 (n_238, in_2[14], n_86);
  nand g195 (out_0[15], n_236, n_237, n_238);
  xor g196 (n_239, in_0[15], in_1[15]);
  xor g197 (n_92, n_239, in_3[15]);
  nand g198 (n_240, in_0[15], in_1[15]);
  nand g199 (n_241, in_3[15], in_1[15]);
  nand g200 (n_242, in_0[15], in_3[15]);
  nand g201 (out_0[16], n_240, n_241, n_242);
  xor g202 (n_243, in_2[15], n_91);
  xor g203 (out_1[15], n_243, n_92);
  nand g204 (n_244, in_2[15], n_91);
  nand g205 (n_245, n_92, n_91);
  nand g206 (n_246, in_2[15], n_92);
  nand g207 (out_1[16], n_244, n_245, n_246);
endmodule

module csa_tree_112_GENERIC(in_0, in_1, in_2, in_3, out_0, out_1);
  input [15:0] in_0, in_1, in_2, in_3;
  output [16:0] out_0, out_1;
  wire [15:0] in_0, in_1, in_2, in_3;
  wire [16:0] out_0, out_1;
  csa_tree_112_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .in_3 (in_3), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_145_229_GENERIC_REAL(in_0, in_1, in_2, in_3, out_0,
     out_1, out_2);
// synthesis_equation "assign out_0 = ( ( in_2 + in_3 ) + ( in_0 * in_1 )  )  ; assign out_1 = 17'b0; assign out_2 = 1'b0;"
  input [15:0] in_0, in_1;
  input [16:0] in_2, in_3;
  output [16:0] out_0, out_1;
  output out_2;
  wire [15:0] in_0, in_1;
  wire [16:0] in_2, in_3;
  wire [16:0] out_0, out_1;
  wire out_2;
  wire n_6, n_8, n_9, n_14, n_15, n_16, n_18, n_19;
  wire n_20, n_22, n_23, n_24, n_26, n_27, n_28, n_30;
  wire n_31, n_32, n_34, n_35, n_36, n_38, n_39, n_40;
  wire n_42, n_43, n_44, n_46, n_47, n_48, n_50, n_51;
  wire n_52, n_54, n_55, n_56, n_58, n_59, n_60, n_62;
  wire n_63, n_64, n_66, n_67, n_68, n_70, n_71, n_72;
  wire n_74, n_75, n_83, n_85, n_86, n_87, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_134, n_136, n_137, n_140, n_142, n_143, n_144, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_185, n_187, n_188, n_191, n_193;
  wire n_194, n_195, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_230, n_232, n_233, n_236, n_238, n_239, n_240, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_269;
  wire n_271, n_272, n_275, n_277, n_278, n_279, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_302, n_304, n_305, n_308, n_310, n_311, n_312, n_316;
  wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_329, n_331, n_332, n_335, n_337;
  wire n_338, n_339, n_343, n_344, n_345, n_346, n_347, n_348;
  wire n_350, n_352, n_353, n_364, n_367, n_368, n_369, n_372;
  wire n_373, n_374, n_375, n_376, n_377, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_476;
  wire n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492;
  wire n_493, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_564;
  wire n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572;
  wire n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580;
  wire n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697;
  wire n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  wire n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761;
  wire n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785;
  wire n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
  wire n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817;
  wire n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841;
  wire n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865;
  wire n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929;
  wire n_930, n_934, n_938, n_942, n_946, n_950, n_954, n_958;
  wire n_962, n_968, n_969, n_970, n_971, n_972, n_973, n_974;
  assign out_2 = in_2[0];
  assign out_0[0] = in_3[0];
  xor g2 (n_6, in_1[1], in_1[0]);
  xor g8 (n_8, in_1[1], in_0[0]);
  and g12 (out_1[0], in_0[0], in_1[0]);
  xor g13 (n_14, in_1[1], in_0[1]);
  nand g14 (n_15, n_14, in_1[0]);
  nand g15 (n_16, n_8, n_9);
  nand g16 (out_0[1], n_15, n_16);
  xor g17 (n_18, in_1[1], in_0[2]);
  nand g18 (n_19, n_18, in_1[0]);
  nand g19 (n_20, n_14, n_9);
  nand g20 (n_369, n_19, n_20);
  xor g21 (n_22, in_1[1], in_0[3]);
  nand g22 (n_23, n_22, in_1[0]);
  nand g23 (n_24, n_18, n_9);
  nand g24 (n_376, n_23, n_24);
  xor g25 (n_26, in_1[1], in_0[4]);
  nand g26 (n_27, n_26, in_1[0]);
  nand g27 (n_28, n_22, n_9);
  nand g28 (n_384, n_27, n_28);
  xor g29 (n_30, in_1[1], in_0[5]);
  nand g30 (n_31, n_30, in_1[0]);
  nand g31 (n_32, n_26, n_9);
  nand g32 (n_394, n_31, n_32);
  xor g33 (n_34, in_1[1], in_0[6]);
  nand g34 (n_35, n_34, in_1[0]);
  nand g35 (n_36, n_30, n_9);
  nand g36 (n_405, n_35, n_36);
  xor g37 (n_38, in_1[1], in_0[7]);
  nand g38 (n_39, n_38, in_1[0]);
  nand g39 (n_40, n_34, n_9);
  nand g40 (n_417, n_39, n_40);
  xor g41 (n_42, in_1[1], in_0[8]);
  nand g42 (n_43, n_42, in_1[0]);
  nand g43 (n_44, n_38, n_9);
  nand g44 (n_432, n_43, n_44);
  xor g45 (n_46, in_1[1], in_0[9]);
  nand g46 (n_47, n_46, in_1[0]);
  nand g47 (n_48, n_42, n_9);
  nand g48 (n_447, n_47, n_48);
  xor g49 (n_50, in_1[1], in_0[10]);
  nand g50 (n_51, n_50, in_1[0]);
  nand g51 (n_52, n_46, n_9);
  nand g52 (n_463, n_51, n_52);
  xor g53 (n_54, in_1[1], in_0[11]);
  nand g54 (n_55, n_54, in_1[0]);
  nand g55 (n_56, n_50, n_9);
  nand g56 (n_484, n_55, n_56);
  xor g57 (n_58, in_1[1], in_0[12]);
  nand g58 (n_59, n_58, in_1[0]);
  nand g59 (n_60, n_54, n_9);
  nand g60 (n_502, n_59, n_60);
  xor g61 (n_62, in_1[1], in_0[13]);
  nand g62 (n_63, n_62, in_1[0]);
  nand g63 (n_64, n_58, n_9);
  nand g64 (n_524, n_63, n_64);
  xor g65 (n_66, in_1[1], in_0[14]);
  nand g66 (n_67, n_66, in_1[0]);
  nand g67 (n_68, n_62, n_9);
  nand g68 (n_547, n_67, n_68);
  xor g69 (n_70, in_1[1], in_0[15]);
  nand g70 (n_71, n_70, in_1[0]);
  nand g71 (n_72, n_66, n_9);
  nand g72 (n_571, n_71, n_72);
  nand g74 (n_74, in_1[1], in_1[0]);
  nand g75 (n_75, n_70, n_9);
  nand g76 (n_598, n_74, n_75);
  xor g81 (n_83, in_1[2], in_1[1]);
  xor g82 (n_85, in_1[3], in_1[2]);
  nor g86 (n_136, in_1[1], in_1[2]);
  nand g87 (n_134, in_1[1], in_1[2]);
  xor g88 (n_86, in_1[3], in_0[0]);
  and g92 (n_368, in_0[0], n_83);
  xor g93 (n_91, in_1[3], in_0[1]);
  nand g94 (n_92, n_91, n_83);
  nand g95 (n_93, n_86, n_87);
  nand g96 (n_375, n_92, n_93);
  xor g97 (n_94, in_1[3], in_0[2]);
  nand g98 (n_95, n_94, n_83);
  nand g99 (n_96, n_91, n_87);
  nand g100 (n_383, n_95, n_96);
  xor g101 (n_97, in_1[3], in_0[3]);
  nand g102 (n_98, n_97, n_83);
  nand g103 (n_99, n_94, n_87);
  nand g104 (n_392, n_98, n_99);
  xor g105 (n_100, in_1[3], in_0[4]);
  nand g106 (n_101, n_100, n_83);
  nand g107 (n_102, n_97, n_87);
  nand g108 (n_402, n_101, n_102);
  xor g109 (n_103, in_1[3], in_0[5]);
  nand g110 (n_104, n_103, n_83);
  nand g111 (n_105, n_100, n_87);
  nand g112 (n_416, n_104, n_105);
  xor g113 (n_106, in_1[3], in_0[6]);
  nand g114 (n_107, n_106, n_83);
  nand g115 (n_108, n_103, n_87);
  nand g116 (n_429, n_107, n_108);
  xor g117 (n_109, in_1[3], in_0[7]);
  nand g118 (n_110, n_109, n_83);
  nand g119 (n_111, n_106, n_87);
  nand g120 (n_443, n_110, n_111);
  xor g121 (n_112, in_1[3], in_0[8]);
  nand g122 (n_113, n_112, n_83);
  nand g123 (n_114, n_109, n_87);
  nand g124 (n_461, n_113, n_114);
  xor g125 (n_115, in_1[3], in_0[9]);
  nand g126 (n_116, n_115, n_83);
  nand g127 (n_117, n_112, n_87);
  nand g128 (n_479, n_116, n_117);
  xor g129 (n_118, in_1[3], in_0[10]);
  nand g130 (n_119, n_118, n_83);
  nand g131 (n_120, n_115, n_87);
  nand g132 (n_500, n_119, n_120);
  xor g133 (n_121, in_1[3], in_0[11]);
  nand g134 (n_122, n_121, n_83);
  nand g135 (n_123, n_118, n_87);
  nand g136 (n_519, n_122, n_123);
  xor g137 (n_124, in_1[3], in_0[12]);
  nand g138 (n_125, n_124, n_83);
  nand g139 (n_126, n_121, n_87);
  nand g140 (n_542, n_125, n_126);
  xor g141 (n_127, in_1[3], in_0[13]);
  nand g142 (n_128, n_127, n_83);
  nand g143 (n_129, n_124, n_87);
  nand g144 (n_567, n_128, n_129);
  xor g145 (n_130, in_1[3], in_0[14]);
  nand g146 (n_131, n_130, n_83);
  nand g147 (n_132, n_127, n_87);
  nand g148 (n_593, n_131, n_132);
  or g151 (n_137, n_968, n_136);
  and g152 (n_374, in_1[3], n_137);
  xor g153 (n_140, in_1[4], in_1[3]);
  xor g154 (n_142, in_1[5], in_1[4]);
  nor g158 (n_187, in_1[3], in_1[4]);
  nand g159 (n_185, in_1[3], in_1[4]);
  xor g160 (n_143, in_1[5], in_0[0]);
  and g164 (n_381, in_0[0], n_140);
  xor g165 (n_148, in_1[5], in_0[1]);
  nand g166 (n_149, n_148, n_140);
  nand g167 (n_150, n_143, n_144);
  nand g168 (n_393, n_149, n_150);
  xor g169 (n_151, in_1[5], in_0[2]);
  nand g170 (n_152, n_151, n_140);
  nand g171 (n_153, n_148, n_144);
  nand g172 (n_404, n_152, n_153);
  xor g173 (n_154, in_1[5], in_0[3]);
  nand g174 (n_155, n_154, n_140);
  nand g175 (n_156, n_151, n_144);
  nand g176 (n_414, n_155, n_156);
  xor g177 (n_157, in_1[5], in_0[4]);
  nand g178 (n_158, n_157, n_140);
  nand g179 (n_159, n_154, n_144);
  nand g180 (n_430, n_158, n_159);
  xor g181 (n_160, in_1[5], in_0[5]);
  nand g182 (n_161, n_160, n_140);
  nand g183 (n_162, n_157, n_144);
  nand g184 (n_445, n_161, n_162);
  xor g185 (n_163, in_1[5], in_0[6]);
  nand g186 (n_164, n_163, n_140);
  nand g187 (n_165, n_160, n_144);
  nand g188 (n_462, n_164, n_165);
  xor g189 (n_166, in_1[5], in_0[7]);
  nand g190 (n_167, n_166, n_140);
  nand g191 (n_168, n_163, n_144);
  nand g192 (n_480, n_167, n_168);
  xor g193 (n_169, in_1[5], in_0[8]);
  nand g194 (n_170, n_169, n_140);
  nand g195 (n_171, n_166, n_144);
  nand g196 (n_501, n_170, n_171);
  xor g197 (n_172, in_1[5], in_0[9]);
  nand g198 (n_173, n_172, n_140);
  nand g199 (n_174, n_169, n_144);
  nand g200 (n_522, n_173, n_174);
  xor g201 (n_175, in_1[5], in_0[10]);
  nand g202 (n_176, n_175, n_140);
  nand g203 (n_177, n_172, n_144);
  nand g204 (n_546, n_176, n_177);
  xor g205 (n_178, in_1[5], in_0[11]);
  nand g206 (n_179, n_178, n_140);
  nand g207 (n_180, n_175, n_144);
  nand g208 (n_570, n_179, n_180);
  xor g209 (n_181, in_1[5], in_0[12]);
  nand g210 (n_182, n_181, n_140);
  nand g211 (n_183, n_178, n_144);
  nand g212 (n_597, n_182, n_183);
  or g215 (n_188, n_969, n_187);
  and g216 (n_390, in_1[5], n_188);
  xor g217 (n_191, in_1[6], in_1[5]);
  xor g218 (n_193, in_1[7], in_1[6]);
  nor g222 (n_232, in_1[5], in_1[6]);
  nand g223 (n_230, in_1[5], in_1[6]);
  xor g224 (n_194, in_1[7], in_0[0]);
  and g228 (n_401, in_0[0], n_191);
  xor g229 (n_199, in_1[7], in_0[1]);
  nand g230 (n_200, n_199, n_191);
  nand g231 (n_201, n_194, n_195);
  nand g232 (n_418, n_200, n_201);
  xor g233 (n_202, in_1[7], in_0[2]);
  nand g234 (n_203, n_202, n_191);
  nand g235 (n_204, n_199, n_195);
  nand g236 (n_431, n_203, n_204);
  xor g237 (n_205, in_1[7], in_0[3]);
  nand g238 (n_206, n_205, n_191);
  nand g239 (n_207, n_202, n_195);
  nand g240 (n_446, n_206, n_207);
  xor g241 (n_208, in_1[7], in_0[4]);
  nand g242 (n_209, n_208, n_191);
  nand g243 (n_210, n_205, n_195);
  nand g244 (n_464, n_209, n_210);
  xor g245 (n_211, in_1[7], in_0[5]);
  nand g246 (n_212, n_211, n_191);
  nand g247 (n_213, n_208, n_195);
  nand g248 (n_483, n_212, n_213);
  xor g249 (n_214, in_1[7], in_0[6]);
  nand g250 (n_215, n_214, n_191);
  nand g251 (n_216, n_211, n_195);
  nand g252 (n_503, n_215, n_216);
  xor g253 (n_217, in_1[7], in_0[7]);
  nand g254 (n_218, n_217, n_191);
  nand g255 (n_219, n_214, n_195);
  nand g256 (n_525, n_218, n_219);
  xor g257 (n_220, in_1[7], in_0[8]);
  nand g258 (n_221, n_220, n_191);
  nand g259 (n_222, n_217, n_195);
  nand g260 (n_548, n_221, n_222);
  xor g261 (n_223, in_1[7], in_0[9]);
  nand g262 (n_224, n_223, n_191);
  nand g263 (n_225, n_220, n_195);
  nand g264 (n_572, n_224, n_225);
  xor g265 (n_226, in_1[7], in_0[10]);
  nand g266 (n_227, n_226, n_191);
  nand g267 (n_228, n_223, n_195);
  nand g268 (n_599, n_227, n_228);
  or g271 (n_233, n_970, n_232);
  and g272 (n_413, in_1[7], n_233);
  xor g273 (n_236, in_1[8], in_1[7]);
  xor g274 (n_238, in_1[9], in_1[8]);
  nor g278 (n_271, in_1[7], in_1[8]);
  nand g279 (n_269, in_1[7], in_1[8]);
  xor g280 (n_239, in_1[9], in_0[0]);
  and g284 (n_427, in_0[0], n_236);
  xor g285 (n_244, in_1[9], in_0[1]);
  nand g286 (n_245, n_244, n_236);
  nand g287 (n_246, n_239, n_240);
  nand g288 (n_448, n_245, n_246);
  xor g289 (n_247, in_1[9], in_0[2]);
  nand g290 (n_248, n_247, n_236);
  nand g291 (n_249, n_244, n_240);
  nand g292 (n_465, n_248, n_249);
  xor g293 (n_250, in_1[9], in_0[3]);
  nand g294 (n_251, n_250, n_236);
  nand g295 (n_252, n_247, n_240);
  nand g296 (n_482, n_251, n_252);
  xor g297 (n_253, in_1[9], in_0[4]);
  nand g298 (n_254, n_253, n_236);
  nand g299 (n_255, n_250, n_240);
  nand g300 (n_504, n_254, n_255);
  xor g301 (n_256, in_1[9], in_0[5]);
  nand g302 (n_257, n_256, n_236);
  nand g303 (n_258, n_253, n_240);
  nand g304 (n_526, n_257, n_258);
  xor g305 (n_259, in_1[9], in_0[6]);
  nand g306 (n_260, n_259, n_236);
  nand g307 (n_261, n_256, n_240);
  nand g308 (n_549, n_260, n_261);
  xor g309 (n_262, in_1[9], in_0[7]);
  nand g310 (n_263, n_262, n_236);
  nand g311 (n_264, n_259, n_240);
  nand g312 (n_574, n_263, n_264);
  xor g313 (n_265, in_1[9], in_0[8]);
  nand g314 (n_266, n_265, n_236);
  nand g315 (n_267, n_262, n_240);
  nand g316 (n_600, n_266, n_267);
  or g319 (n_272, n_971, n_271);
  and g320 (n_442, in_1[9], n_272);
  xor g321 (n_275, in_1[10], in_1[9]);
  xor g322 (n_277, in_1[11], in_1[10]);
  nor g326 (n_304, in_1[9], in_1[10]);
  nand g327 (n_302, in_1[9], in_1[10]);
  xor g328 (n_278, in_1[11], in_0[0]);
  and g332 (n_459, in_0[0], n_275);
  xor g333 (n_283, in_1[11], in_0[1]);
  nand g334 (n_284, n_283, n_275);
  nand g335 (n_285, n_278, n_279);
  nand g336 (n_478, n_284, n_285);
  xor g337 (n_286, in_1[11], in_0[2]);
  nand g338 (n_287, n_286, n_275);
  nand g339 (n_288, n_283, n_279);
  nand g340 (n_499, n_287, n_288);
  xor g341 (n_289, in_1[11], in_0[3]);
  nand g342 (n_290, n_289, n_275);
  nand g343 (n_291, n_286, n_279);
  nand g344 (n_520, n_290, n_291);
  xor g345 (n_292, in_1[11], in_0[4]);
  nand g346 (n_293, n_292, n_275);
  nand g347 (n_294, n_289, n_279);
  nand g348 (n_543, n_293, n_294);
  xor g349 (n_295, in_1[11], in_0[5]);
  nand g350 (n_296, n_295, n_275);
  nand g351 (n_297, n_292, n_279);
  nand g352 (n_568, n_296, n_297);
  xor g353 (n_298, in_1[11], in_0[6]);
  nand g354 (n_299, n_298, n_275);
  nand g355 (n_300, n_295, n_279);
  nand g356 (n_594, n_299, n_300);
  or g359 (n_305, n_972, n_304);
  and g360 (n_477, in_1[11], n_305);
  xor g361 (n_308, in_1[12], in_1[11]);
  xor g362 (n_310, in_1[13], in_1[12]);
  nor g366 (n_331, in_1[11], in_1[12]);
  nand g367 (n_329, in_1[11], in_1[12]);
  xor g368 (n_311, in_1[13], in_0[0]);
  and g372 (n_497, in_0[0], n_308);
  xor g373 (n_316, in_1[13], in_0[1]);
  nand g374 (n_317, n_316, n_308);
  nand g375 (n_318, n_311, n_312);
  nand g376 (n_521, n_317, n_318);
  xor g377 (n_319, in_1[13], in_0[2]);
  nand g378 (n_320, n_319, n_308);
  nand g379 (n_321, n_316, n_312);
  nand g380 (n_545, n_320, n_321);
  xor g381 (n_322, in_1[13], in_0[3]);
  nand g382 (n_323, n_322, n_308);
  nand g383 (n_324, n_319, n_312);
  nand g384 (n_566, n_323, n_324);
  xor g385 (n_325, in_1[13], in_0[4]);
  nand g386 (n_326, n_325, n_308);
  nand g387 (n_327, n_322, n_312);
  nand g388 (n_595, n_326, n_327);
  or g391 (n_332, n_973, n_331);
  and g392 (n_518, in_1[13], n_332);
  xor g393 (n_335, in_1[14], in_1[13]);
  xor g394 (n_337, in_1[15], in_1[14]);
  nor g398 (n_352, in_1[13], in_1[14]);
  nand g399 (n_350, in_1[13], in_1[14]);
  xor g400 (n_338, in_1[15], in_0[0]);
  and g404 (n_541, in_0[0], n_335);
  xor g405 (n_343, in_1[15], in_0[1]);
  nand g406 (n_344, n_343, n_335);
  nand g407 (n_345, n_338, n_339);
  nand g408 (n_569, n_344, n_345);
  xor g409 (n_346, in_1[15], in_0[2]);
  nand g410 (n_347, n_346, n_335);
  nand g411 (n_348, n_343, n_339);
  nand g412 (n_596, n_347, n_348);
  or g415 (n_353, n_974, n_352);
  and g416 (n_565, in_1[15], n_353);
  and g428 (n_591, in_0[0], in_1[15]);
  xor g516 (n_650, in_2[1], in_3[1]);
  xor g517 (out_1[1], n_650, n_364);
  nand g518 (n_651, in_2[1], in_3[1]);
  nand g519 (n_652, n_364, in_3[1]);
  nand g520 (n_653, in_2[1], n_364);
  nand g521 (out_0[2], n_651, n_652, n_653);
  xor g522 (n_367, in_2[2], in_3[2]);
  and g523 (n_372, in_2[2], in_3[2]);
  xor g524 (n_654, n_367, n_368);
  xor g525 (out_1[2], n_654, n_369);
  nand g526 (n_655, n_367, n_368);
  nand g527 (n_656, n_369, n_368);
  nand g528 (n_657, n_367, n_369);
  nand g529 (out_0[3], n_655, n_656, n_657);
  xor g530 (n_373, in_2[3], in_3[3]);
  and g531 (n_380, in_2[3], in_3[3]);
  xor g532 (n_658, n_372, n_373);
  xor g533 (n_377, n_658, n_374);
  nand g534 (n_659, n_372, n_373);
  nand g535 (n_660, n_374, n_373);
  nand g536 (n_661, n_372, n_374);
  nand g537 (n_385, n_659, n_660, n_661);
  xor g538 (n_662, n_375, n_376);
  xor g539 (out_1[3], n_662, n_377);
  nand g540 (n_663, n_375, n_376);
  nand g541 (n_664, n_377, n_376);
  nand g542 (n_665, n_375, n_377);
  nand g543 (n_386, n_663, n_664, n_665);
  xor g544 (n_666, in_2[4], in_3[4]);
  xor g545 (n_382, n_666, n_380);
  nand g546 (n_667, in_2[4], in_3[4]);
  nand g547 (n_668, n_380, in_3[4]);
  nand g548 (n_669, in_2[4], n_380);
  nand g549 (n_391, n_667, n_668, n_669);
  xor g550 (n_670, n_381, n_382);
  xor g551 (out_0[4], n_670, n_383);
  nand g552 (n_671, n_381, n_382);
  nand g553 (n_672, n_383, n_382);
  nand g554 (n_673, n_381, n_383);
  nand g555 (n_395, n_671, n_672, n_673);
  xor g556 (n_674, n_384, n_385);
  xor g557 (out_1[4], n_674, n_386);
  nand g558 (n_675, n_384, n_385);
  nand g559 (n_676, n_386, n_385);
  nand g560 (n_677, n_384, n_386);
  nand g561 (out_0[5], n_675, n_676, n_677);
  xor g562 (n_389, in_2[5], in_3[5]);
  and g563 (n_400, in_2[5], in_3[5]);
  xor g564 (n_678, n_389, n_390);
  xor g565 (n_396, n_678, n_391);
  nand g566 (n_679, n_389, n_390);
  nand g567 (n_680, n_391, n_390);
  nand g568 (n_681, n_389, n_391);
  nand g569 (n_407, n_679, n_680, n_681);
  xor g570 (n_682, n_392, n_393);
  xor g571 (n_397, n_682, n_394);
  nand g572 (n_683, n_392, n_393);
  nand g573 (n_684, n_394, n_393);
  nand g574 (n_685, n_392, n_394);
  nand g575 (n_406, n_683, n_684, n_685);
  xor g576 (n_686, n_395, n_396);
  xor g577 (out_1[5], n_686, n_397);
  nand g578 (n_687, n_395, n_396);
  nand g579 (n_688, n_397, n_396);
  nand g580 (n_689, n_395, n_397);
  nand g581 (out_0[6], n_687, n_688, n_689);
  xor g582 (n_690, in_2[6], in_3[6]);
  xor g583 (n_403, n_690, n_400);
  nand g584 (n_691, in_2[6], in_3[6]);
  nand g585 (n_692, n_400, in_3[6]);
  nand g586 (n_693, in_2[6], n_400);
  nand g587 (n_415, n_691, n_692, n_693);
  xor g588 (n_694, n_401, n_402);
  xor g589 (n_408, n_694, n_403);
  nand g590 (n_695, n_401, n_402);
  nand g591 (n_696, n_403, n_402);
  nand g592 (n_697, n_401, n_403);
  nand g593 (n_420, n_695, n_696, n_697);
  xor g594 (n_698, n_404, n_405);
  xor g595 (n_409, n_698, n_406);
  nand g596 (n_699, n_404, n_405);
  nand g597 (n_700, n_406, n_405);
  nand g598 (n_701, n_404, n_406);
  nand g599 (n_422, n_699, n_700, n_701);
  xor g600 (n_702, n_407, n_408);
  xor g601 (out_1[6], n_702, n_409);
  nand g602 (n_703, n_407, n_408);
  nand g603 (n_704, n_409, n_408);
  nand g604 (n_705, n_407, n_409);
  nand g605 (out_0[7], n_703, n_704, n_705);
  xor g606 (n_412, in_2[7], in_3[7]);
  and g607 (n_426, in_2[7], in_3[7]);
  xor g608 (n_706, n_412, n_413);
  xor g609 (n_419, n_706, n_414);
  nand g610 (n_707, n_412, n_413);
  nand g611 (n_708, n_414, n_413);
  nand g612 (n_709, n_412, n_414);
  nand g613 (n_433, n_707, n_708, n_709);
  xor g614 (n_710, n_415, n_416);
  xor g615 (n_421, n_710, n_417);
  nand g616 (n_711, n_415, n_416);
  nand g617 (n_712, n_417, n_416);
  nand g618 (n_713, n_415, n_417);
  nand g619 (n_434, n_711, n_712, n_713);
  xor g620 (n_714, n_418, n_419);
  xor g621 (n_423, n_714, n_420);
  nand g622 (n_715, n_418, n_419);
  nand g623 (n_716, n_420, n_419);
  nand g624 (n_717, n_418, n_420);
  nand g625 (n_437, n_715, n_716, n_717);
  xor g626 (n_718, n_421, n_422);
  xor g627 (out_1[7], n_718, n_423);
  nand g628 (n_719, n_421, n_422);
  nand g629 (n_720, n_423, n_422);
  nand g630 (n_721, n_421, n_423);
  nand g631 (out_0[8], n_719, n_720, n_721);
  xor g632 (n_722, in_2[8], in_3[8]);
  xor g633 (n_428, n_722, n_426);
  nand g634 (n_723, in_2[8], in_3[8]);
  nand g635 (n_724, n_426, in_3[8]);
  nand g636 (n_725, in_2[8], n_426);
  nand g637 (n_444, n_723, n_724, n_725);
  xor g638 (n_726, n_427, n_428);
  xor g639 (n_435, n_726, n_429);
  nand g640 (n_727, n_427, n_428);
  nand g641 (n_728, n_429, n_428);
  nand g642 (n_729, n_427, n_429);
  nand g643 (n_451, n_727, n_728, n_729);
  xor g644 (n_730, n_430, n_431);
  xor g645 (n_436, n_730, n_432);
  nand g646 (n_731, n_430, n_431);
  nand g647 (n_732, n_432, n_431);
  nand g648 (n_733, n_430, n_432);
  nand g649 (n_450, n_731, n_732, n_733);
  xor g650 (n_734, n_433, n_434);
  xor g651 (n_438, n_734, n_435);
  nand g652 (n_735, n_433, n_434);
  nand g653 (n_736, n_435, n_434);
  nand g654 (n_737, n_433, n_435);
  nand g655 (n_455, n_735, n_736, n_737);
  xor g656 (n_738, n_436, n_437);
  xor g657 (out_1[8], n_738, n_438);
  nand g658 (n_739, n_436, n_437);
  nand g659 (n_740, n_438, n_437);
  nand g660 (n_741, n_436, n_438);
  nand g661 (out_0[9], n_739, n_740, n_741);
  xor g662 (n_441, in_2[9], in_3[9]);
  and g663 (n_458, in_2[9], in_3[9]);
  xor g664 (n_742, n_441, n_442);
  xor g665 (n_449, n_742, n_443);
  nand g666 (n_743, n_441, n_442);
  nand g667 (n_744, n_443, n_442);
  nand g668 (n_745, n_441, n_443);
  nand g669 (n_466, n_743, n_744, n_745);
  xor g670 (n_746, n_444, n_445);
  xor g671 (n_452, n_746, n_446);
  nand g672 (n_747, n_444, n_445);
  nand g673 (n_748, n_446, n_445);
  nand g674 (n_749, n_444, n_446);
  nand g675 (n_467, n_747, n_748, n_749);
  xor g676 (n_750, n_447, n_448);
  xor g677 (n_453, n_750, n_449);
  nand g678 (n_751, n_447, n_448);
  nand g679 (n_752, n_449, n_448);
  nand g680 (n_753, n_447, n_449);
  nand g681 (n_470, n_751, n_752, n_753);
  xor g682 (n_754, n_450, n_451);
  xor g683 (n_454, n_754, n_452);
  nand g684 (n_755, n_450, n_451);
  nand g685 (n_756, n_452, n_451);
  nand g686 (n_757, n_450, n_452);
  nand g687 (n_471, n_755, n_756, n_757);
  xor g688 (n_758, n_453, n_454);
  xor g689 (out_1[9], n_758, n_455);
  nand g690 (n_759, n_453, n_454);
  nand g691 (n_760, n_455, n_454);
  nand g692 (n_761, n_453, n_455);
  nand g693 (out_0[10], n_759, n_760, n_761);
  xor g694 (n_762, in_2[10], in_3[10]);
  xor g695 (n_460, n_762, n_458);
  nand g696 (n_763, in_2[10], in_3[10]);
  nand g697 (n_764, n_458, in_3[10]);
  nand g698 (n_765, in_2[10], n_458);
  nand g699 (n_481, n_763, n_764, n_765);
  xor g700 (n_766, n_459, n_460);
  xor g701 (n_469, n_766, n_461);
  nand g702 (n_767, n_459, n_460);
  nand g703 (n_768, n_461, n_460);
  nand g704 (n_769, n_459, n_461);
  nand g705 (n_485, n_767, n_768, n_769);
  xor g706 (n_770, n_462, n_463);
  xor g707 (n_468, n_770, n_464);
  nand g708 (n_771, n_462, n_463);
  nand g709 (n_772, n_464, n_463);
  nand g710 (n_773, n_462, n_464);
  nand g711 (n_487, n_771, n_772, n_773);
  xor g712 (n_774, n_465, n_466);
  xor g713 (n_472, n_774, n_467);
  nand g714 (n_775, n_465, n_466);
  nand g715 (n_776, n_467, n_466);
  nand g716 (n_777, n_465, n_467);
  nand g717 (n_490, n_775, n_776, n_777);
  xor g718 (n_778, n_468, n_469);
  xor g719 (n_473, n_778, n_470);
  nand g720 (n_779, n_468, n_469);
  nand g721 (n_780, n_470, n_469);
  nand g722 (n_781, n_468, n_470);
  nand g723 (n_493, n_779, n_780, n_781);
  xor g724 (n_782, n_471, n_472);
  xor g725 (out_1[10], n_782, n_473);
  nand g726 (n_783, n_471, n_472);
  nand g727 (n_784, n_473, n_472);
  nand g728 (n_785, n_471, n_473);
  nand g729 (out_0[11], n_783, n_784, n_785);
  xor g730 (n_476, in_2[11], in_3[11]);
  and g731 (n_496, in_2[11], in_3[11]);
  xor g732 (n_786, n_476, n_477);
  xor g733 (n_486, n_786, n_478);
  nand g734 (n_787, n_476, n_477);
  nand g735 (n_788, n_478, n_477);
  nand g736 (n_789, n_476, n_478);
  nand g737 (n_507, n_787, n_788, n_789);
  xor g738 (n_790, n_479, n_480);
  xor g739 (n_489, n_790, n_481);
  nand g740 (n_791, n_479, n_480);
  nand g741 (n_792, n_481, n_480);
  nand g742 (n_793, n_479, n_481);
  nand g743 (n_506, n_791, n_792, n_793);
  xor g744 (n_794, n_482, n_483);
  xor g745 (n_488, n_794, n_484);
  nand g746 (n_795, n_482, n_483);
  nand g747 (n_796, n_484, n_483);
  nand g748 (n_797, n_482, n_484);
  nand g749 (n_505, n_795, n_796, n_797);
  xor g750 (n_798, n_485, n_486);
  xor g751 (n_491, n_798, n_487);
  nand g752 (n_799, n_485, n_486);
  nand g753 (n_800, n_487, n_486);
  nand g754 (n_801, n_485, n_487);
  nand g755 (n_511, n_799, n_800, n_801);
  xor g756 (n_802, n_488, n_489);
  xor g757 (n_492, n_802, n_490);
  nand g758 (n_803, n_488, n_489);
  nand g759 (n_804, n_490, n_489);
  nand g760 (n_805, n_488, n_490);
  nand g761 (n_513, n_803, n_804, n_805);
  xor g762 (n_806, n_491, n_492);
  xor g763 (out_1[11], n_806, n_493);
  nand g764 (n_807, n_491, n_492);
  nand g765 (n_808, n_493, n_492);
  nand g766 (n_809, n_491, n_493);
  nand g767 (out_0[12], n_807, n_808, n_809);
  xor g768 (n_810, in_2[12], in_3[12]);
  xor g769 (n_498, n_810, n_496);
  nand g770 (n_811, in_2[12], in_3[12]);
  nand g771 (n_812, n_496, in_3[12]);
  nand g772 (n_813, in_2[12], n_496);
  nand g773 (n_523, n_811, n_812, n_813);
  xor g774 (n_814, n_497, n_498);
  xor g775 (n_508, n_814, n_499);
  nand g776 (n_815, n_497, n_498);
  nand g777 (n_816, n_499, n_498);
  nand g778 (n_817, n_497, n_499);
  nand g779 (n_527, n_815, n_816, n_817);
  xor g780 (n_818, n_500, n_501);
  xor g781 (n_509, n_818, n_502);
  nand g782 (n_819, n_500, n_501);
  nand g783 (n_820, n_502, n_501);
  nand g784 (n_821, n_500, n_502);
  nand g785 (n_528, n_819, n_820, n_821);
  xor g786 (n_822, n_503, n_504);
  xor g787 (n_510, n_822, n_505);
  nand g788 (n_823, n_503, n_504);
  nand g789 (n_824, n_505, n_504);
  nand g790 (n_825, n_503, n_505);
  nand g791 (n_532, n_823, n_824, n_825);
  xor g792 (n_826, n_506, n_507);
  xor g793 (n_512, n_826, n_508);
  nand g794 (n_827, n_506, n_507);
  nand g795 (n_828, n_508, n_507);
  nand g796 (n_829, n_506, n_508);
  nand g797 (n_534, n_827, n_828, n_829);
  xor g798 (n_830, n_509, n_510);
  xor g799 (n_514, n_830, n_511);
  nand g800 (n_831, n_509, n_510);
  nand g801 (n_832, n_511, n_510);
  nand g802 (n_833, n_509, n_511);
  nand g803 (n_536, n_831, n_832, n_833);
  xor g804 (n_834, n_512, n_513);
  xor g805 (out_1[12], n_834, n_514);
  nand g806 (n_835, n_512, n_513);
  nand g807 (n_836, n_514, n_513);
  nand g808 (n_837, n_512, n_514);
  nand g809 (out_0[13], n_835, n_836, n_837);
  xor g810 (n_517, in_2[13], in_3[13]);
  and g811 (n_540, in_2[13], in_3[13]);
  xor g812 (n_838, n_517, n_518);
  xor g813 (n_529, n_838, n_519);
  nand g814 (n_839, n_517, n_518);
  nand g815 (n_840, n_519, n_518);
  nand g816 (n_841, n_517, n_519);
  nand g817 (n_552, n_839, n_840, n_841);
  xor g818 (n_842, n_520, n_521);
  xor g819 (n_531, n_842, n_522);
  nand g820 (n_843, n_520, n_521);
  nand g821 (n_844, n_522, n_521);
  nand g822 (n_845, n_520, n_522);
  nand g823 (n_550, n_843, n_844, n_845);
  xor g824 (n_846, n_523, n_524);
  xor g825 (n_530, n_846, n_525);
  nand g826 (n_847, n_523, n_524);
  nand g827 (n_848, n_525, n_524);
  nand g828 (n_849, n_523, n_525);
  nand g829 (n_551, n_847, n_848, n_849);
  xor g830 (n_850, n_526, n_527);
  xor g831 (n_533, n_850, n_528);
  nand g832 (n_851, n_526, n_527);
  nand g833 (n_852, n_528, n_527);
  nand g834 (n_853, n_526, n_528);
  nand g835 (n_556, n_851, n_852, n_853);
  xor g836 (n_854, n_529, n_530);
  xor g837 (n_535, n_854, n_531);
  nand g838 (n_855, n_529, n_530);
  nand g839 (n_856, n_531, n_530);
  nand g840 (n_857, n_529, n_531);
  nand g841 (n_558, n_855, n_856, n_857);
  xor g842 (n_858, n_532, n_533);
  xor g843 (n_537, n_858, n_534);
  nand g844 (n_859, n_532, n_533);
  nand g845 (n_860, n_534, n_533);
  nand g846 (n_861, n_532, n_534);
  nand g847 (n_560, n_859, n_860, n_861);
  xor g848 (n_862, n_535, n_536);
  xor g849 (out_1[13], n_862, n_537);
  nand g850 (n_863, n_535, n_536);
  nand g851 (n_864, n_537, n_536);
  nand g852 (n_865, n_535, n_537);
  nand g853 (out_0[14], n_863, n_864, n_865);
  xor g854 (n_866, in_2[14], in_3[14]);
  xor g855 (n_544, n_866, n_540);
  nand g856 (n_867, in_2[14], in_3[14]);
  nand g857 (n_868, n_540, in_3[14]);
  nand g858 (n_869, in_2[14], n_540);
  nand g859 (n_573, n_867, n_868, n_869);
  xor g860 (n_870, n_541, n_542);
  xor g861 (n_554, n_870, n_543);
  nand g862 (n_871, n_541, n_542);
  nand g863 (n_872, n_543, n_542);
  nand g864 (n_873, n_541, n_543);
  nand g865 (n_578, n_871, n_872, n_873);
  xor g866 (n_874, n_544, n_545);
  xor g867 (n_555, n_874, n_546);
  nand g868 (n_875, n_544, n_545);
  nand g869 (n_876, n_546, n_545);
  nand g870 (n_877, n_544, n_546);
  nand g871 (n_575, n_875, n_876, n_877);
  xor g872 (n_878, n_547, n_548);
  xor g873 (n_553, n_878, n_549);
  nand g874 (n_879, n_547, n_548);
  nand g875 (n_880, n_549, n_548);
  nand g876 (n_881, n_547, n_549);
  nand g877 (n_577, n_879, n_880, n_881);
  xor g878 (n_882, n_550, n_551);
  xor g879 (n_557, n_882, n_552);
  nand g880 (n_883, n_550, n_551);
  nand g881 (n_884, n_552, n_551);
  nand g882 (n_885, n_550, n_552);
  nand g883 (n_581, n_883, n_884, n_885);
  xor g884 (n_886, n_553, n_554);
  xor g885 (n_559, n_886, n_555);
  nand g886 (n_887, n_553, n_554);
  nand g887 (n_888, n_555, n_554);
  nand g888 (n_889, n_553, n_555);
  nand g889 (n_583, n_887, n_888, n_889);
  xor g890 (n_890, n_556, n_557);
  xor g891 (n_561, n_890, n_558);
  nand g892 (n_891, n_556, n_557);
  nand g893 (n_892, n_558, n_557);
  nand g894 (n_893, n_556, n_558);
  nand g895 (n_586, n_891, n_892, n_893);
  xor g896 (n_894, n_559, n_560);
  xor g897 (out_1[14], n_894, n_561);
  nand g898 (n_895, n_559, n_560);
  nand g899 (n_896, n_561, n_560);
  nand g900 (n_897, n_559, n_561);
  nand g901 (out_0[15], n_895, n_896, n_897);
  xor g902 (n_564, in_2[15], in_3[15]);
  and g903 (n_590, in_2[15], in_3[15]);
  xor g904 (n_898, n_564, n_565);
  xor g905 (n_576, n_898, n_566);
  nand g906 (n_899, n_564, n_565);
  nand g907 (n_900, n_566, n_565);
  nand g908 (n_901, n_564, n_566);
  nand g909 (n_603, n_899, n_900, n_901);
  xor g910 (n_902, n_567, n_568);
  xor g911 (n_580, n_902, n_569);
  nand g912 (n_903, n_567, n_568);
  nand g913 (n_904, n_569, n_568);
  nand g914 (n_905, n_567, n_569);
  nand g915 (n_601, n_903, n_904, n_905);
  xor g916 (n_906, n_570, n_571);
  xor g917 (n_579, n_906, n_572);
  nand g918 (n_907, n_570, n_571);
  nand g919 (n_908, n_572, n_571);
  nand g920 (n_909, n_570, n_572);
  nand g921 (n_602, n_907, n_908, n_909);
  xor g922 (n_910, n_573, n_574);
  xor g923 (n_582, n_910, n_575);
  nand g924 (n_911, n_573, n_574);
  nand g925 (n_912, n_575, n_574);
  nand g926 (n_913, n_573, n_575);
  nand g927 (n_607, n_911, n_912, n_913);
  xor g928 (n_914, n_576, n_577);
  xor g929 (n_584, n_914, n_578);
  nand g930 (n_915, n_576, n_577);
  nand g931 (n_916, n_578, n_577);
  nand g932 (n_917, n_576, n_578);
  nand g933 (n_608, n_915, n_916, n_917);
  xor g934 (n_918, n_579, n_580);
  xor g935 (n_585, n_918, n_581);
  nand g936 (n_919, n_579, n_580);
  nand g937 (n_920, n_581, n_580);
  nand g938 (n_921, n_579, n_581);
  nand g939 (n_611, n_919, n_920, n_921);
  xor g940 (n_922, n_582, n_583);
  xor g941 (n_587, n_922, n_584);
  nand g942 (n_923, n_582, n_583);
  nand g943 (n_924, n_584, n_583);
  nand g944 (n_925, n_582, n_584);
  nand g945 (n_613, n_923, n_924, n_925);
  xor g946 (n_926, n_585, n_586);
  xor g947 (out_1[15], n_926, n_587);
  nand g948 (n_927, n_585, n_586);
  nand g949 (n_928, n_587, n_586);
  nand g950 (n_929, n_585, n_587);
  nand g951 (out_0[16], n_927, n_928, n_929);
  xor g952 (n_930, in_2[16], in_3[16]);
  xor g953 (n_592, n_930, n_590);
  xor g958 (n_934, n_591, n_592);
  xor g959 (n_604, n_934, n_593);
  xor g964 (n_938, n_594, n_595);
  xor g965 (n_606, n_938, n_596);
  xor g970 (n_942, n_597, n_598);
  xor g971 (n_605, n_942, n_599);
  xor g976 (n_946, n_600, n_601);
  xor g977 (n_609, n_946, n_602);
  xor g982 (n_950, n_603, n_604);
  xor g983 (n_610, n_950, n_605);
  xor g988 (n_954, n_606, n_607);
  xor g989 (n_612, n_954, n_608);
  xor g994 (n_958, n_609, n_610);
  xor g995 (n_614, n_958, n_611);
  xor g1000 (n_962, n_612, n_613);
  xor g1001 (out_1[16], n_962, n_614);
  and g1007 (n_968, wc, n_134);
  not gc (wc, in_0[0]);
  and g1008 (n_969, wc0, n_185);
  not gc0 (wc0, in_0[0]);
  and g1009 (n_970, wc1, n_230);
  not gc1 (wc1, in_0[0]);
  and g1010 (n_971, wc2, n_269);
  not gc2 (wc2, in_0[0]);
  and g1011 (n_972, wc3, n_302);
  not gc3 (wc3, in_0[0]);
  and g1012 (n_973, wc4, n_329);
  not gc4 (wc4, in_0[0]);
  and g1013 (n_974, wc5, n_350);
  not gc5 (wc5, in_0[0]);
  and g1014 (n_9, wc6, n_6);
  not gc6 (wc6, in_1[0]);
  and g1016 (n_87, n_85, wc7);
  not gc7 (wc7, n_83);
  and g1017 (n_144, n_142, wc8);
  not gc8 (wc8, n_140);
  and g1018 (n_195, n_193, wc9);
  not gc9 (wc9, n_191);
  and g1019 (n_240, n_238, wc10);
  not gc10 (wc10, n_236);
  and g1020 (n_279, n_277, wc11);
  not gc11 (wc11, n_275);
  and g1021 (n_312, n_310, wc12);
  not gc12 (wc12, n_308);
  and g1022 (n_339, n_337, wc13);
  not gc13 (wc13, n_335);
  and g1023 (n_364, in_1[1], wc14);
  not gc14 (wc14, out_1[0]);
endmodule

module csa_tree_145_229_GENERIC(in_0, in_1, in_2, in_3, out_0, out_1,
     out_2);
  input [15:0] in_0, in_1;
  input [16:0] in_2, in_3;
  output [16:0] out_0, out_1;
  output out_2;
  wire [15:0] in_0, in_1;
  wire [16:0] in_2, in_3;
  wire [16:0] out_0, out_1;
  wire out_2;
  csa_tree_145_229_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .in_3 (in_3), .out_0 (out_0), .out_1 (out_1), .out_2
       (out_2));
endmodule

module csa_tree_31_GENERIC_REAL(in_0, in_1, out_0, out_1);
// synthesis_equation "assign out_0 = ( in_0 * in_1 )  ; assign out_1 = 16'b0;"
  input [7:0] in_0, in_1;
  output [15:0] out_0, out_1;
  wire [7:0] in_0, in_1;
  wire [15:0] out_0, out_1;
  wire n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305;
  assign out_1[0] = 1'b0;
  assign out_1[15] = 1'b0;
  assign out_0[15] = 1'b0;
  and g1 (out_0[0], in_0[0], in_1[0]);
  and g2 (out_0[1], in_0[1], in_1[0]);
  and g3 (n_17, in_0[2], in_1[0]);
  and g4 (n_19, in_0[3], in_1[0]);
  and g5 (n_24, in_0[4], in_1[0]);
  and g6 (n_32, in_0[5], in_1[0]);
  and g7 (n_43, in_0[6], in_1[0]);
  and g8 (n_57, in_0[7], in_1[0]);
  and g9 (out_1[1], in_0[0], in_1[1]);
  and g10 (out_0[2], in_0[1], in_1[1]);
  and g11 (n_20, in_0[2], in_1[1]);
  and g12 (n_25, in_0[3], in_1[1]);
  and g13 (n_33, in_0[4], in_1[1]);
  and g14 (n_44, in_0[5], in_1[1]);
  and g15 (n_58, in_0[6], in_1[1]);
  and g16 (n_74, in_0[7], in_1[1]);
  and g17 (n_18, in_0[0], in_1[2]);
  and g18 (n_22, in_0[1], in_1[2]);
  and g19 (n_28, in_0[2], in_1[2]);
  and g20 (n_36, in_0[3], in_1[2]);
  and g21 (n_47, in_0[4], in_1[2]);
  and g22 (n_62, in_0[5], in_1[2]);
  and g23 (n_75, in_0[6], in_1[2]);
  and g24 (n_91, in_0[7], in_1[2]);
  and g25 (n_21, in_0[0], in_1[3]);
  and g26 (n_26, in_0[1], in_1[3]);
  and g27 (n_34, in_0[2], in_1[3]);
  and g28 (n_45, in_0[3], in_1[3]);
  and g29 (n_59, in_0[4], in_1[3]);
  and g30 (n_78, in_0[5], in_1[3]);
  and g31 (n_92, in_0[6], in_1[3]);
  and g32 (n_106, in_0[7], in_1[3]);
  and g33 (n_27, in_0[0], in_1[4]);
  and g34 (n_35, in_0[1], in_1[4]);
  and g35 (n_46, in_0[2], in_1[4]);
  and g36 (n_61, in_0[3], in_1[4]);
  and g37 (n_76, in_0[4], in_1[4]);
  and g38 (n_95, in_0[5], in_1[4]);
  and g39 (n_107, in_0[6], in_1[4]);
  and g40 (n_118, in_0[7], in_1[4]);
  and g41 (n_37, in_0[0], in_1[5]);
  and g42 (n_48, in_0[1], in_1[5]);
  and g43 (n_63, in_0[2], in_1[5]);
  and g44 (n_77, in_0[3], in_1[5]);
  and g45 (n_93, in_0[4], in_1[5]);
  and g46 (n_110, in_0[5], in_1[5]);
  and g47 (n_119, in_0[6], in_1[5]);
  and g48 (n_127, in_0[7], in_1[5]);
  and g49 (n_49, in_0[0], in_1[6]);
  and g50 (n_64, in_0[1], in_1[6]);
  and g51 (n_79, in_0[2], in_1[6]);
  and g52 (n_94, in_0[3], in_1[6]);
  and g53 (n_108, in_0[4], in_1[6]);
  and g54 (n_121, in_0[5], in_1[6]);
  and g55 (n_128, in_0[6], in_1[6]);
  and g56 (n_133, in_0[7], in_1[6]);
  and g57 (n_60, in_0[0], in_1[7]);
  and g58 (n_80, in_0[1], in_1[7]);
  and g59 (n_96, in_0[2], in_1[7]);
  and g60 (n_109, in_0[3], in_1[7]);
  and g61 (n_120, in_0[4], in_1[7]);
  and g62 (n_129, in_0[5], in_1[7]);
  and g63 (n_134, in_0[6], in_1[7]);
  and g64 (out_0[14], in_0[7], in_1[7]);
  xor g107 (out_1[2], n_17, n_18);
  and g108 (out_0[3], n_17, n_18);
  xor g109 (n_23, n_19, n_20);
  and g110 (n_30, n_19, n_20);
  xor g111 (n_166, n_21, n_22);
  xor g112 (out_1[3], n_166, n_23);
  nand g113 (n_167, n_21, n_22);
  nand g114 (n_168, n_23, n_22);
  nand g115 (n_169, n_21, n_23);
  nand g116 (out_0[4], n_167, n_168, n_169);
  xor g117 (n_29, n_24, n_25);
  and g118 (n_39, n_24, n_25);
  xor g119 (n_170, n_26, n_27);
  xor g120 (n_31, n_170, n_28);
  nand g121 (n_171, n_26, n_27);
  nand g122 (n_172, n_28, n_27);
  nand g123 (n_173, n_26, n_28);
  nand g124 (n_40, n_171, n_172, n_173);
  xor g125 (n_174, n_29, n_30);
  xor g126 (out_1[4], n_174, n_31);
  nand g127 (n_175, n_29, n_30);
  nand g128 (n_176, n_31, n_30);
  nand g129 (n_177, n_29, n_31);
  nand g130 (out_0[5], n_175, n_176, n_177);
  xor g131 (n_38, n_32, n_33);
  and g132 (n_50, n_32, n_33);
  xor g133 (n_178, n_34, n_35);
  xor g134 (n_41, n_178, n_36);
  nand g135 (n_179, n_34, n_35);
  nand g136 (n_180, n_36, n_35);
  nand g137 (n_181, n_34, n_36);
  nand g138 (n_52, n_179, n_180, n_181);
  xor g139 (n_182, n_37, n_38);
  xor g140 (n_42, n_182, n_39);
  nand g141 (n_183, n_37, n_38);
  nand g142 (n_184, n_39, n_38);
  nand g143 (n_185, n_37, n_39);
  nand g144 (n_54, n_183, n_184, n_185);
  xor g145 (n_186, n_40, n_41);
  xor g146 (out_1[5], n_186, n_42);
  nand g147 (n_187, n_40, n_41);
  nand g148 (n_188, n_42, n_41);
  nand g149 (n_189, n_40, n_42);
  nand g150 (out_0[6], n_187, n_188, n_189);
  xor g151 (n_51, n_43, n_44);
  and g152 (n_65, n_43, n_44);
  xor g153 (n_190, n_45, n_46);
  xor g154 (n_53, n_190, n_47);
  nand g155 (n_191, n_45, n_46);
  nand g156 (n_192, n_47, n_46);
  nand g157 (n_193, n_45, n_47);
  nand g158 (n_67, n_191, n_192, n_193);
  xor g159 (n_194, n_48, n_49);
  xor g160 (n_55, n_194, n_50);
  nand g161 (n_195, n_48, n_49);
  nand g162 (n_196, n_50, n_49);
  nand g163 (n_197, n_48, n_50);
  nand g164 (n_70, n_195, n_196, n_197);
  xor g165 (n_198, n_51, n_52);
  xor g166 (n_56, n_198, n_53);
  nand g167 (n_199, n_51, n_52);
  nand g168 (n_200, n_53, n_52);
  nand g169 (n_201, n_51, n_53);
  nand g170 (n_72, n_199, n_200, n_201);
  xor g171 (n_202, n_54, n_55);
  xor g172 (out_1[6], n_202, n_56);
  nand g173 (n_203, n_54, n_55);
  nand g174 (n_204, n_56, n_55);
  nand g175 (n_205, n_54, n_56);
  nand g176 (out_0[7], n_203, n_204, n_205);
  xor g177 (n_66, n_57, n_58);
  and g178 (n_82, n_57, n_58);
  xor g179 (n_206, n_59, n_60);
  xor g180 (n_69, n_206, n_61);
  nand g181 (n_207, n_59, n_60);
  nand g182 (n_208, n_61, n_60);
  nand g183 (n_209, n_59, n_61);
  nand g184 (n_83, n_207, n_208, n_209);
  xor g185 (n_210, n_62, n_63);
  xor g186 (n_68, n_210, n_64);
  nand g187 (n_211, n_62, n_63);
  nand g188 (n_212, n_64, n_63);
  nand g189 (n_213, n_62, n_64);
  nand g190 (n_84, n_211, n_212, n_213);
  xor g191 (n_214, n_65, n_66);
  xor g192 (n_71, n_214, n_67);
  nand g193 (n_215, n_65, n_66);
  nand g194 (n_216, n_67, n_66);
  nand g195 (n_217, n_65, n_67);
  nand g196 (n_87, n_215, n_216, n_217);
  xor g197 (n_218, n_68, n_69);
  xor g198 (n_73, n_218, n_70);
  nand g199 (n_219, n_68, n_69);
  nand g200 (n_220, n_70, n_69);
  nand g201 (n_221, n_68, n_70);
  nand g202 (n_89, n_219, n_220, n_221);
  xor g203 (n_222, n_71, n_72);
  xor g204 (out_1[7], n_222, n_73);
  nand g205 (n_223, n_71, n_72);
  nand g206 (n_224, n_73, n_72);
  nand g207 (n_225, n_71, n_73);
  nand g208 (out_0[8], n_223, n_224, n_225);
  xor g209 (n_81, n_74, n_75);
  and g210 (n_97, n_74, n_75);
  xor g211 (n_226, n_76, n_77);
  xor g212 (n_85, n_226, n_78);
  nand g213 (n_227, n_76, n_77);
  nand g214 (n_228, n_78, n_77);
  nand g215 (n_229, n_76, n_78);
  nand g216 (n_98, n_227, n_228, n_229);
  xor g217 (n_230, n_79, n_80);
  xor g218 (n_86, n_230, n_81);
  nand g219 (n_231, n_79, n_80);
  nand g220 (n_232, n_81, n_80);
  nand g221 (n_233, n_79, n_81);
  nand g222 (n_101, n_231, n_232, n_233);
  xor g223 (n_234, n_82, n_83);
  xor g224 (n_88, n_234, n_84);
  nand g225 (n_235, n_82, n_83);
  nand g226 (n_236, n_84, n_83);
  nand g227 (n_237, n_82, n_84);
  nand g228 (n_102, n_235, n_236, n_237);
  xor g229 (n_238, n_85, n_86);
  xor g230 (n_90, n_238, n_87);
  nand g231 (n_239, n_85, n_86);
  nand g232 (n_240, n_87, n_86);
  nand g233 (n_241, n_85, n_87);
  nand g234 (n_105, n_239, n_240, n_241);
  xor g235 (n_242, n_88, n_89);
  xor g236 (out_1[8], n_242, n_90);
  nand g237 (n_243, n_88, n_89);
  nand g238 (n_244, n_90, n_89);
  nand g239 (n_245, n_88, n_90);
  nand g240 (out_0[9], n_243, n_244, n_245);
  xor g241 (n_246, n_91, n_92);
  xor g242 (n_100, n_246, n_93);
  nand g243 (n_247, n_91, n_92);
  nand g244 (n_248, n_93, n_92);
  nand g245 (n_249, n_91, n_93);
  nand g246 (n_112, n_247, n_248, n_249);
  xor g247 (n_250, n_94, n_95);
  xor g248 (n_99, n_250, n_96);
  nand g249 (n_251, n_94, n_95);
  nand g250 (n_252, n_96, n_95);
  nand g251 (n_253, n_94, n_96);
  nand g252 (n_111, n_251, n_252, n_253);
  xor g253 (n_254, n_97, n_98);
  xor g254 (n_103, n_254, n_99);
  nand g255 (n_255, n_97, n_98);
  nand g256 (n_256, n_99, n_98);
  nand g257 (n_257, n_97, n_99);
  nand g258 (n_115, n_255, n_256, n_257);
  xor g259 (n_258, n_100, n_101);
  xor g260 (n_104, n_258, n_102);
  nand g261 (n_259, n_100, n_101);
  nand g262 (n_260, n_102, n_101);
  nand g263 (n_261, n_100, n_102);
  nand g264 (n_117, n_259, n_260, n_261);
  xor g265 (n_262, n_103, n_104);
  xor g266 (out_1[9], n_262, n_105);
  nand g267 (n_263, n_103, n_104);
  nand g268 (n_264, n_105, n_104);
  nand g269 (n_265, n_103, n_105);
  nand g270 (out_0[10], n_263, n_264, n_265);
  xor g271 (n_266, n_106, n_107);
  xor g272 (n_113, n_266, n_108);
  nand g273 (n_267, n_106, n_107);
  nand g274 (n_268, n_108, n_107);
  nand g275 (n_269, n_106, n_108);
  nand g276 (n_122, n_267, n_268, n_269);
  xor g277 (n_270, n_109, n_110);
  xor g278 (n_114, n_270, n_111);
  nand g279 (n_271, n_109, n_110);
  nand g280 (n_272, n_111, n_110);
  nand g281 (n_273, n_109, n_111);
  nand g282 (n_124, n_271, n_272, n_273);
  xor g283 (n_274, n_112, n_113);
  xor g284 (n_116, n_274, n_114);
  nand g285 (n_275, n_112, n_113);
  nand g286 (n_276, n_114, n_113);
  nand g287 (n_277, n_112, n_114);
  nand g288 (n_126, n_275, n_276, n_277);
  xor g289 (n_278, n_115, n_116);
  xor g290 (out_1[10], n_278, n_117);
  nand g291 (n_279, n_115, n_116);
  nand g292 (n_280, n_117, n_116);
  nand g293 (n_281, n_115, n_117);
  nand g294 (out_0[11], n_279, n_280, n_281);
  xor g295 (n_282, n_118, n_119);
  xor g296 (n_123, n_282, n_120);
  nand g297 (n_283, n_118, n_119);
  nand g298 (n_284, n_120, n_119);
  nand g299 (n_285, n_118, n_120);
  nand g300 (n_130, n_283, n_284, n_285);
  xor g301 (n_286, n_121, n_122);
  xor g302 (n_125, n_286, n_123);
  nand g303 (n_287, n_121, n_122);
  nand g304 (n_288, n_123, n_122);
  nand g305 (n_289, n_121, n_123);
  nand g306 (n_132, n_287, n_288, n_289);
  xor g307 (n_290, n_124, n_125);
  xor g308 (out_1[11], n_290, n_126);
  nand g309 (n_291, n_124, n_125);
  nand g310 (n_292, n_126, n_125);
  nand g311 (n_293, n_124, n_126);
  nand g312 (out_1[12], n_291, n_292, n_293);
  xor g313 (n_294, n_127, n_128);
  xor g314 (n_131, n_294, n_129);
  nand g315 (n_295, n_127, n_128);
  nand g316 (n_296, n_129, n_128);
  nand g317 (n_297, n_127, n_129);
  nand g318 (n_135, n_295, n_296, n_297);
  xor g319 (n_298, n_130, n_131);
  xor g320 (out_0[12], n_298, n_132);
  nand g321 (n_299, n_130, n_131);
  nand g322 (n_300, n_132, n_131);
  nand g323 (n_301, n_130, n_132);
  nand g324 (out_1[13], n_299, n_300, n_301);
  xor g325 (n_302, n_133, n_134);
  xor g326 (out_0[13], n_302, n_135);
  nand g327 (n_303, n_133, n_134);
  nand g328 (n_304, n_135, n_134);
  nand g329 (n_305, n_133, n_135);
  nand g330 (out_1[14], n_303, n_304, n_305);
endmodule

module csa_tree_31_GENERIC(in_0, in_1, out_0, out_1);
  input [7:0] in_0, in_1;
  output [15:0] out_0, out_1;
  wire [7:0] in_0, in_1;
  wire [15:0] out_0, out_1;
  csa_tree_31_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .out_0
       (out_0), .out_1 (out_1));
endmodule

