library verilog;
use verilog.vl_types.all;
entity Distance_tb is
end Distance_tb;
