library verilog;
use verilog.vl_types.all;
entity p2s_tb is
end p2s_tb;
