module csa_tree_add_53_18_group_20_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( in_2 + ( in_0 * in_1 )  )  ;"
  input [7:0] in_0;
  input [3:0] in_1;
  input [9:0] in_2;
  output [9:0] out_0;
  wire [7:0] in_0;
  wire [3:0] in_1;
  wire [9:0] in_2;
  wire [9:0] out_0;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_181, n_186, n_188, n_191, n_193, n_194, n_196, n_198;
  wire n_199, n_201, n_203, n_204, n_206, n_208, n_209, n_211;
  wire n_213, n_214, n_216, n_218, n_219, n_221, n_223, n_224;
  wire n_226, n_228, n_229, n_231, n_243, n_244, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260;
  and g1 (n_42, in_0[0], in_1[0]);
  and g2 (n_41, in_0[1], in_1[0]);
  and g3 (n_55, in_0[2], in_1[0]);
  and g4 (n_59, in_0[3], in_1[0]);
  and g5 (n_66, in_0[4], in_1[0]);
  and g6 (n_74, in_0[5], in_1[0]);
  and g7 (n_82, in_0[6], in_1[0]);
  and g8 (n_89, in_0[7], in_1[0]);
  and g9 (n_54, in_0[0], in_1[1]);
  and g10 (n_57, in_0[1], in_1[1]);
  and g11 (n_62, in_0[2], in_1[1]);
  and g12 (n_69, in_0[3], in_1[1]);
  and g13 (n_77, in_0[4], in_1[1]);
  and g14 (n_85, in_0[5], in_1[1]);
  and g15 (n_92, in_0[6], in_1[1]);
  and g16 (n_97, in_0[7], in_1[1]);
  and g17 (n_56, in_0[0], in_1[2]);
  and g18 (n_60, in_0[1], in_1[2]);
  and g19 (n_67, in_0[2], in_1[2]);
  and g20 (n_75, in_0[3], in_1[2]);
  and g21 (n_83, in_0[4], in_1[2]);
  and g22 (n_90, in_0[5], in_1[2]);
  and g23 (n_99, in_0[6], in_1[2]);
  and g24 (n_104, in_0[7], in_1[2]);
  and g25 (n_61, in_0[0], in_1[3]);
  and g26 (n_68, in_0[1], in_1[3]);
  and g27 (n_76, in_0[2], in_1[3]);
  and g28 (n_84, in_0[3], in_1[3]);
  and g29 (n_91, in_0[4], in_1[3]);
  and g30 (n_98, in_0[5], in_1[3]);
  and g31 (n_105, in_0[6], in_1[3]);
  xor g55 (n_51, in_2[1], n_54);
  and g56 (n_40, in_2[1], n_54);
  xor g57 (n_58, in_2[2], n_55);
  and g58 (n_64, in_2[2], n_55);
  xor g59 (n_109, n_56, n_57);
  xor g60 (n_50, n_109, n_58);
  nand g61 (n_110, n_56, n_57);
  nand g62 (n_111, n_58, n_57);
  nand g63 (n_112, n_56, n_58);
  nand g64 (n_39, n_110, n_111, n_112);
  xor g65 (n_63, in_2[3], n_59);
  and g66 (n_70, in_2[3], n_59);
  xor g67 (n_113, n_60, n_61);
  xor g68 (n_65, n_113, n_62);
  nand g69 (n_114, n_60, n_61);
  nand g70 (n_115, n_62, n_61);
  nand g71 (n_116, n_60, n_62);
  nand g72 (n_71, n_114, n_115, n_116);
  xor g73 (n_117, n_63, n_64);
  xor g74 (n_49, n_117, n_65);
  nand g75 (n_118, n_63, n_64);
  nand g76 (n_119, n_65, n_64);
  nand g77 (n_120, n_63, n_65);
  nand g78 (n_38, n_118, n_119, n_120);
  xor g79 (n_121, in_2[4], n_66);
  xor g80 (n_72, n_121, n_67);
  nand g81 (n_122, in_2[4], n_66);
  nand g82 (n_123, n_67, n_66);
  nand g83 (n_124, in_2[4], n_67);
  nand g84 (n_78, n_122, n_123, n_124);
  xor g85 (n_125, n_68, n_69);
  xor g86 (n_73, n_125, n_70);
  nand g87 (n_126, n_68, n_69);
  nand g88 (n_127, n_70, n_69);
  nand g89 (n_128, n_68, n_70);
  nand g90 (n_80, n_126, n_127, n_128);
  xor g91 (n_129, n_71, n_72);
  xor g92 (n_48, n_129, n_73);
  nand g93 (n_130, n_71, n_72);
  nand g94 (n_131, n_73, n_72);
  nand g95 (n_132, n_71, n_73);
  nand g96 (n_37, n_130, n_131, n_132);
  xor g97 (n_133, in_2[5], n_74);
  xor g98 (n_79, n_133, n_75);
  nand g99 (n_134, in_2[5], n_74);
  nand g100 (n_135, n_75, n_74);
  nand g101 (n_136, in_2[5], n_75);
  nand g102 (n_86, n_134, n_135, n_136);
  xor g103 (n_137, n_76, n_77);
  xor g104 (n_81, n_137, n_78);
  nand g105 (n_138, n_76, n_77);
  nand g106 (n_139, n_78, n_77);
  nand g107 (n_140, n_76, n_78);
  nand g108 (n_88, n_138, n_139, n_140);
  xor g109 (n_141, n_79, n_80);
  xor g110 (n_47, n_141, n_81);
  nand g111 (n_142, n_79, n_80);
  nand g112 (n_143, n_81, n_80);
  nand g113 (n_144, n_79, n_81);
  nand g114 (n_36, n_142, n_143, n_144);
  xor g115 (n_145, in_2[6], n_82);
  xor g116 (n_87, n_145, n_83);
  nand g117 (n_146, in_2[6], n_82);
  nand g118 (n_147, n_83, n_82);
  nand g119 (n_148, in_2[6], n_83);
  nand g120 (n_93, n_146, n_147, n_148);
  xor g121 (n_149, n_84, n_85);
  xor g122 (n_53, n_149, n_86);
  nand g123 (n_150, n_84, n_85);
  nand g124 (n_151, n_86, n_85);
  nand g125 (n_152, n_84, n_86);
  nand g126 (n_96, n_150, n_151, n_152);
  xor g127 (n_153, n_87, n_53);
  xor g128 (n_46, n_153, n_88);
  nand g129 (n_154, n_87, n_53);
  nand g130 (n_155, n_88, n_53);
  nand g131 (n_156, n_87, n_88);
  nand g132 (n_35, n_154, n_155, n_156);
  xor g133 (n_157, in_2[7], n_89);
  xor g134 (n_94, n_157, n_90);
  nand g135 (n_158, in_2[7], n_89);
  nand g136 (n_159, n_90, n_89);
  nand g137 (n_160, in_2[7], n_90);
  nand g138 (n_101, n_158, n_159, n_160);
  xor g139 (n_161, n_91, n_92);
  xor g140 (n_95, n_161, n_93);
  nand g141 (n_162, n_91, n_92);
  nand g142 (n_163, n_93, n_92);
  nand g143 (n_164, n_91, n_93);
  nand g144 (n_103, n_162, n_163, n_164);
  xor g145 (n_165, n_94, n_95);
  xor g146 (n_45, n_165, n_96);
  nand g147 (n_166, n_94, n_95);
  nand g148 (n_167, n_96, n_95);
  nand g149 (n_168, n_94, n_96);
  nand g150 (n_34, n_166, n_167, n_168);
  xor g151 (n_100, in_2[8], n_97);
  and g152 (n_106, in_2[8], n_97);
  xor g153 (n_169, n_98, n_99);
  xor g154 (n_102, n_169, n_100);
  nand g155 (n_170, n_98, n_99);
  nand g156 (n_171, n_100, n_99);
  nand g157 (n_172, n_98, n_100);
  nand g158 (n_108, n_170, n_171, n_172);
  xor g159 (n_173, n_101, n_102);
  xor g160 (n_44, n_173, n_103);
  nand g161 (n_174, n_101, n_102);
  nand g162 (n_175, n_103, n_102);
  nand g163 (n_176, n_101, n_103);
  nand g164 (n_43, n_174, n_175, n_176);
  xor g165 (n_177, in_2[9], n_104);
  xor g166 (n_107, n_177, n_105);
  xor g171 (n_181, n_106, n_107);
  xor g172 (n_33, n_181, n_108);
  nand g179 (n_186, n_42, in_2[0]);
  nor g182 (n_188, n_41, n_51);
  nand g183 (n_191, n_41, n_51);
  nor g184 (n_193, n_40, n_50);
  nand g185 (n_196, n_40, n_50);
  nor g186 (n_198, n_39, n_49);
  nand g187 (n_201, n_39, n_49);
  nor g188 (n_203, n_38, n_48);
  nand g189 (n_206, n_38, n_48);
  nor g190 (n_208, n_37, n_47);
  nand g191 (n_211, n_37, n_47);
  nor g192 (n_213, n_36, n_46);
  nand g193 (n_216, n_36, n_46);
  nor g194 (n_218, n_35, n_45);
  nand g195 (n_221, n_35, n_45);
  nor g196 (n_223, n_34, n_44);
  nand g197 (n_226, n_34, n_44);
  nor g198 (n_228, n_33, n_43);
  nand g199 (n_231, n_33, n_43);
  nand g202 (n_194, n_191, n_243);
  nand g205 (n_199, n_196, n_247);
  nand g32 (n_204, n_201, n_250);
  nand g35 (n_209, n_206, n_256);
  nand g38 (n_214, n_211, n_257);
  nand g41 (n_219, n_216, n_258);
  nand g44 (n_224, n_221, n_259);
  nand g47 (n_229, n_226, n_260);
  xnor g54 (out_0[2], n_194, n_246);
  xnor g209 (out_0[3], n_199, n_248);
  xnor g211 (out_0[4], n_204, n_249);
  xnor g213 (out_0[5], n_209, n_251);
  xnor g215 (out_0[6], n_214, n_252);
  xnor g217 (out_0[7], n_219, n_253);
  xnor g219 (out_0[8], n_224, n_254);
  xnor g221 (out_0[9], n_229, n_255);
  xor g222 (out_0[0], in_2[0], n_42);
  or g224 (n_243, n_186, n_188);
  or g225 (n_244, wc, n_188);
  not gc (wc, n_191);
  xor g226 (out_0[1], n_186, n_244);
  or g227 (n_246, wc0, n_193);
  not gc0 (wc0, n_196);
  or g228 (n_247, wc1, n_193);
  not gc1 (wc1, n_194);
  or g229 (n_248, wc2, n_198);
  not gc2 (wc2, n_201);
  or g230 (n_249, wc3, n_203);
  not gc3 (wc3, n_206);
  or g231 (n_250, wc4, n_198);
  not gc4 (wc4, n_199);
  or g232 (n_251, wc5, n_208);
  not gc5 (wc5, n_211);
  or g233 (n_252, wc6, n_213);
  not gc6 (wc6, n_216);
  or g234 (n_253, wc7, n_218);
  not gc7 (wc7, n_221);
  or g235 (n_254, wc8, n_223);
  not gc8 (wc8, n_226);
  or g236 (n_255, wc9, n_228);
  not gc9 (wc9, n_231);
  or g237 (n_256, wc10, n_203);
  not gc10 (wc10, n_204);
  or g238 (n_257, wc11, n_208);
  not gc11 (wc11, n_209);
  or g239 (n_258, wc12, n_213);
  not gc12 (wc12, n_214);
  or g240 (n_259, wc13, n_218);
  not gc13 (wc13, n_219);
  or g241 (n_260, wc14, n_223);
  not gc14 (wc14, n_224);
endmodule

module csa_tree_add_53_18_group_20_GENERIC(in_0, in_1, in_2, out_0);
  input [7:0] in_0;
  input [3:0] in_1;
  input [9:0] in_2;
  output [9:0] out_0;
  wire [7:0] in_0;
  wire [3:0] in_1;
  wire [9:0] in_2;
  wire [9:0] out_0;
  csa_tree_add_53_18_group_20_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_54_18_group_22_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( in_2 + ( in_0 * in_1 )  )  ;"
  input [7:0] in_0;
  input [3:0] in_1;
  input [9:0] in_2;
  output [9:0] out_0;
  wire [7:0] in_0;
  wire [3:0] in_1;
  wire [9:0] in_2;
  wire [9:0] out_0;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_181, n_186, n_188, n_191, n_193, n_194, n_196, n_198;
  wire n_199, n_201, n_203, n_204, n_206, n_208, n_209, n_211;
  wire n_213, n_214, n_216, n_218, n_219, n_221, n_223, n_224;
  wire n_226, n_228, n_229, n_231, n_243, n_244, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260;
  and g1 (n_42, in_0[0], in_1[0]);
  and g2 (n_41, in_0[1], in_1[0]);
  and g3 (n_55, in_0[2], in_1[0]);
  and g4 (n_59, in_0[3], in_1[0]);
  and g5 (n_66, in_0[4], in_1[0]);
  and g6 (n_74, in_0[5], in_1[0]);
  and g7 (n_82, in_0[6], in_1[0]);
  and g8 (n_89, in_0[7], in_1[0]);
  and g9 (n_54, in_0[0], in_1[1]);
  and g10 (n_57, in_0[1], in_1[1]);
  and g11 (n_62, in_0[2], in_1[1]);
  and g12 (n_69, in_0[3], in_1[1]);
  and g13 (n_77, in_0[4], in_1[1]);
  and g14 (n_85, in_0[5], in_1[1]);
  and g15 (n_92, in_0[6], in_1[1]);
  and g16 (n_97, in_0[7], in_1[1]);
  and g17 (n_56, in_0[0], in_1[2]);
  and g18 (n_60, in_0[1], in_1[2]);
  and g19 (n_67, in_0[2], in_1[2]);
  and g20 (n_75, in_0[3], in_1[2]);
  and g21 (n_83, in_0[4], in_1[2]);
  and g22 (n_90, in_0[5], in_1[2]);
  and g23 (n_99, in_0[6], in_1[2]);
  and g24 (n_104, in_0[7], in_1[2]);
  and g25 (n_61, in_0[0], in_1[3]);
  and g26 (n_68, in_0[1], in_1[3]);
  and g27 (n_76, in_0[2], in_1[3]);
  and g28 (n_84, in_0[3], in_1[3]);
  and g29 (n_91, in_0[4], in_1[3]);
  and g30 (n_98, in_0[5], in_1[3]);
  and g31 (n_105, in_0[6], in_1[3]);
  xor g55 (n_51, in_2[1], n_54);
  and g56 (n_40, in_2[1], n_54);
  xor g57 (n_58, in_2[2], n_55);
  and g58 (n_64, in_2[2], n_55);
  xor g59 (n_109, n_56, n_57);
  xor g60 (n_50, n_109, n_58);
  nand g61 (n_110, n_56, n_57);
  nand g62 (n_111, n_58, n_57);
  nand g63 (n_112, n_56, n_58);
  nand g64 (n_39, n_110, n_111, n_112);
  xor g65 (n_63, in_2[3], n_59);
  and g66 (n_70, in_2[3], n_59);
  xor g67 (n_113, n_60, n_61);
  xor g68 (n_65, n_113, n_62);
  nand g69 (n_114, n_60, n_61);
  nand g70 (n_115, n_62, n_61);
  nand g71 (n_116, n_60, n_62);
  nand g72 (n_71, n_114, n_115, n_116);
  xor g73 (n_117, n_63, n_64);
  xor g74 (n_49, n_117, n_65);
  nand g75 (n_118, n_63, n_64);
  nand g76 (n_119, n_65, n_64);
  nand g77 (n_120, n_63, n_65);
  nand g78 (n_38, n_118, n_119, n_120);
  xor g79 (n_121, in_2[4], n_66);
  xor g80 (n_72, n_121, n_67);
  nand g81 (n_122, in_2[4], n_66);
  nand g82 (n_123, n_67, n_66);
  nand g83 (n_124, in_2[4], n_67);
  nand g84 (n_78, n_122, n_123, n_124);
  xor g85 (n_125, n_68, n_69);
  xor g86 (n_73, n_125, n_70);
  nand g87 (n_126, n_68, n_69);
  nand g88 (n_127, n_70, n_69);
  nand g89 (n_128, n_68, n_70);
  nand g90 (n_80, n_126, n_127, n_128);
  xor g91 (n_129, n_71, n_72);
  xor g92 (n_48, n_129, n_73);
  nand g93 (n_130, n_71, n_72);
  nand g94 (n_131, n_73, n_72);
  nand g95 (n_132, n_71, n_73);
  nand g96 (n_37, n_130, n_131, n_132);
  xor g97 (n_133, in_2[5], n_74);
  xor g98 (n_79, n_133, n_75);
  nand g99 (n_134, in_2[5], n_74);
  nand g100 (n_135, n_75, n_74);
  nand g101 (n_136, in_2[5], n_75);
  nand g102 (n_86, n_134, n_135, n_136);
  xor g103 (n_137, n_76, n_77);
  xor g104 (n_81, n_137, n_78);
  nand g105 (n_138, n_76, n_77);
  nand g106 (n_139, n_78, n_77);
  nand g107 (n_140, n_76, n_78);
  nand g108 (n_88, n_138, n_139, n_140);
  xor g109 (n_141, n_79, n_80);
  xor g110 (n_47, n_141, n_81);
  nand g111 (n_142, n_79, n_80);
  nand g112 (n_143, n_81, n_80);
  nand g113 (n_144, n_79, n_81);
  nand g114 (n_36, n_142, n_143, n_144);
  xor g115 (n_145, in_2[6], n_82);
  xor g116 (n_87, n_145, n_83);
  nand g117 (n_146, in_2[6], n_82);
  nand g118 (n_147, n_83, n_82);
  nand g119 (n_148, in_2[6], n_83);
  nand g120 (n_93, n_146, n_147, n_148);
  xor g121 (n_149, n_84, n_85);
  xor g122 (n_53, n_149, n_86);
  nand g123 (n_150, n_84, n_85);
  nand g124 (n_151, n_86, n_85);
  nand g125 (n_152, n_84, n_86);
  nand g126 (n_96, n_150, n_151, n_152);
  xor g127 (n_153, n_87, n_53);
  xor g128 (n_46, n_153, n_88);
  nand g129 (n_154, n_87, n_53);
  nand g130 (n_155, n_88, n_53);
  nand g131 (n_156, n_87, n_88);
  nand g132 (n_35, n_154, n_155, n_156);
  xor g133 (n_157, in_2[7], n_89);
  xor g134 (n_94, n_157, n_90);
  nand g135 (n_158, in_2[7], n_89);
  nand g136 (n_159, n_90, n_89);
  nand g137 (n_160, in_2[7], n_90);
  nand g138 (n_101, n_158, n_159, n_160);
  xor g139 (n_161, n_91, n_92);
  xor g140 (n_95, n_161, n_93);
  nand g141 (n_162, n_91, n_92);
  nand g142 (n_163, n_93, n_92);
  nand g143 (n_164, n_91, n_93);
  nand g144 (n_103, n_162, n_163, n_164);
  xor g145 (n_165, n_94, n_95);
  xor g146 (n_45, n_165, n_96);
  nand g147 (n_166, n_94, n_95);
  nand g148 (n_167, n_96, n_95);
  nand g149 (n_168, n_94, n_96);
  nand g150 (n_34, n_166, n_167, n_168);
  xor g151 (n_100, in_2[8], n_97);
  and g152 (n_106, in_2[8], n_97);
  xor g153 (n_169, n_98, n_99);
  xor g154 (n_102, n_169, n_100);
  nand g155 (n_170, n_98, n_99);
  nand g156 (n_171, n_100, n_99);
  nand g157 (n_172, n_98, n_100);
  nand g158 (n_108, n_170, n_171, n_172);
  xor g159 (n_173, n_101, n_102);
  xor g160 (n_44, n_173, n_103);
  nand g161 (n_174, n_101, n_102);
  nand g162 (n_175, n_103, n_102);
  nand g163 (n_176, n_101, n_103);
  nand g164 (n_43, n_174, n_175, n_176);
  xor g165 (n_177, in_2[9], n_104);
  xor g166 (n_107, n_177, n_105);
  xor g171 (n_181, n_106, n_107);
  xor g172 (n_33, n_181, n_108);
  nand g179 (n_186, n_42, in_2[0]);
  nor g182 (n_188, n_41, n_51);
  nand g183 (n_191, n_41, n_51);
  nor g184 (n_193, n_40, n_50);
  nand g185 (n_196, n_40, n_50);
  nor g186 (n_198, n_39, n_49);
  nand g187 (n_201, n_39, n_49);
  nor g188 (n_203, n_38, n_48);
  nand g189 (n_206, n_38, n_48);
  nor g190 (n_208, n_37, n_47);
  nand g191 (n_211, n_37, n_47);
  nor g192 (n_213, n_36, n_46);
  nand g193 (n_216, n_36, n_46);
  nor g194 (n_218, n_35, n_45);
  nand g195 (n_221, n_35, n_45);
  nor g196 (n_223, n_34, n_44);
  nand g197 (n_226, n_34, n_44);
  nor g198 (n_228, n_33, n_43);
  nand g199 (n_231, n_33, n_43);
  nand g202 (n_194, n_191, n_243);
  nand g205 (n_199, n_196, n_247);
  nand g32 (n_204, n_201, n_250);
  nand g35 (n_209, n_206, n_256);
  nand g38 (n_214, n_211, n_257);
  nand g41 (n_219, n_216, n_258);
  nand g44 (n_224, n_221, n_259);
  nand g47 (n_229, n_226, n_260);
  xnor g54 (out_0[2], n_194, n_246);
  xnor g209 (out_0[3], n_199, n_248);
  xnor g211 (out_0[4], n_204, n_249);
  xnor g213 (out_0[5], n_209, n_251);
  xnor g215 (out_0[6], n_214, n_252);
  xnor g217 (out_0[7], n_219, n_253);
  xnor g219 (out_0[8], n_224, n_254);
  xnor g221 (out_0[9], n_229, n_255);
  xor g222 (out_0[0], in_2[0], n_42);
  or g224 (n_243, n_186, n_188);
  or g225 (n_244, wc, n_188);
  not gc (wc, n_191);
  xor g226 (out_0[1], n_186, n_244);
  or g227 (n_246, wc0, n_193);
  not gc0 (wc0, n_196);
  or g228 (n_247, wc1, n_193);
  not gc1 (wc1, n_194);
  or g229 (n_248, wc2, n_198);
  not gc2 (wc2, n_201);
  or g230 (n_249, wc3, n_203);
  not gc3 (wc3, n_206);
  or g231 (n_250, wc4, n_198);
  not gc4 (wc4, n_199);
  or g232 (n_251, wc5, n_208);
  not gc5 (wc5, n_211);
  or g233 (n_252, wc6, n_213);
  not gc6 (wc6, n_216);
  or g234 (n_253, wc7, n_218);
  not gc7 (wc7, n_221);
  or g235 (n_254, wc8, n_223);
  not gc8 (wc8, n_226);
  or g236 (n_255, wc9, n_228);
  not gc9 (wc9, n_231);
  or g237 (n_256, wc10, n_203);
  not gc10 (wc10, n_204);
  or g238 (n_257, wc11, n_208);
  not gc11 (wc11, n_209);
  or g239 (n_258, wc12, n_213);
  not gc12 (wc12, n_214);
  or g240 (n_259, wc13, n_218);
  not gc13 (wc13, n_219);
  or g241 (n_260, wc14, n_223);
  not gc14 (wc14, n_224);
endmodule

module csa_tree_add_54_18_group_22_GENERIC(in_0, in_1, in_2, out_0);
  input [7:0] in_0;
  input [3:0] in_1;
  input [9:0] in_2;
  output [9:0] out_0;
  wire [7:0] in_0;
  wire [3:0] in_1;
  wire [9:0] in_2;
  wire [9:0] out_0;
  csa_tree_add_54_18_group_22_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module divide_unsigned_GENERIC_REAL(A, B, QUOTIENT);
// synthesis_equation "assign QUOTIENT = A / B;"
  input [9:0] A, B;
  output [9:0] QUOTIENT;
  wire [9:0] A, B;
  wire [9:0] QUOTIENT;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_42, n_43, n_44, n_46, n_47, n_49, n_50, n_53;
  wire n_54, n_56, n_57, n_58, n_59, n_60, n_61, n_62;
  wire n_63, n_64, n_66, n_67, n_69, n_70, n_73, n_74;
  wire n_75, n_76, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_94, n_95, n_97, n_98, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_109, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_132, n_133, n_135, n_136, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_186, n_198, n_204, n_206;
  wire n_207, n_208, n_209, n_212, n_213, n_214, n_215, n_218;
  wire n_219, n_220, n_221, n_223, n_224, n_228, n_231, n_233;
  wire n_234, n_235, n_237, n_239, n_244, n_247, n_252, n_256;
  wire n_260, n_264, n_268, n_270, n_273, n_276, n_277, n_282;
  wire n_284, n_286, n_289, n_290, n_291, n_301, n_307, n_318;
  wire n_321, n_323, n_326, n_327, n_340, n_363, n_365, n_368;
  wire n_369, n_370, n_372, n_373, n_375, n_383, n_393, n_410;
  wire n_412, n_414, n_415, n_416, n_417, n_419, n_420, n_423;
  wire n_425, n_429, n_446, n_458, n_461, n_463, n_464, n_465;
  wire n_466, n_468, n_469, n_472, n_474, n_480, n_499, n_515;
  wire n_517, n_518, n_519, n_520, n_522, n_523, n_526, n_528;
  wire n_535, n_557, n_574, n_576, n_578, n_579, n_580, n_581;
  wire n_583, n_584, n_585, n_586, n_587, n_589, n_590, n_593;
  wire n_595, n_598, n_603, n_610, n_620, n_624, n_639, n_642;
  wire n_644, n_645, n_646, n_647, n_649, n_650, n_651, n_652;
  wire n_653, n_655, n_656, n_659, n_661, n_664, n_671, n_678;
  wire n_690, n_694, n_713, n_715, n_716, n_717, n_718, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_727, n_730, n_732;
  wire n_735, n_743, n_750, n_765, n_769, n_789, n_791, n_793;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_802;
  wire n_804, n_805, n_806, n_807, n_808, n_810, n_811, n_814;
  wire n_816, n_817, n_818, n_820, n_822, n_827, n_830, n_835;
  wire n_839, n_846, n_850, n_852, n_855, n_868, n_871, n_873;
  wire n_874, n_875, n_876, n_878, n_879, n_880, n_881, n_882;
  wire n_884, n_885, n_886, n_887, n_888, n_890, n_891, n_894;
  wire n_896, n_897, n_898, n_900, n_902, n_909, n_912, n_917;
  wire n_921, n_930, n_934, n_936, n_939, n_956, n_958, n_959;
  wire n_960, n_961, n_963, n_964, n_965, n_966, n_967, n_969;
  wire n_970, n_971, n_972, n_973, n_975, n_976, n_979, n_981;
  wire n_982, n_983, n_985, n_987, n_995, n_998, n_1003, n_1007;
  wire n_1019, n_1023, n_1025, n_1028, n_1045, n_1047, n_1052, n_1054;
  wire n_1058, n_1060, n_1064, n_1066, n_1070, n_1072, n_1075, n_1078;
  wire n_1080, n_1084, n_1086, n_1091, n_1099, n_1103, n_1106, n_1108;
  wire n_1146, n_1148, n_1152, n_1154, n_1158, n_1160, n_1164, n_1166;
  wire n_1169, n_1172, n_1174, n_1178, n_1180, n_1186, n_1187, n_1189;
  wire n_1197, n_1201, n_1247, n_1249, n_1253, n_1255, n_1259, n_1261;
  wire n_1265, n_1267, n_1270, n_1273, n_1275, n_1279, n_1281, n_1288;
  wire n_1293, n_1301, n_1305, n_1312, n_1342, n_1343, n_1344, n_1345;
  wire n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353;
  wire n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361;
  wire n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369;
  wire n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377;
  wire n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385;
  wire n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393;
  wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
  wire n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409;
  wire n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418;
  wire n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1427;
  wire n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435;
  wire n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443;
  wire n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468;
  wire n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484;
  wire n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508;
  wire n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517;
  wire n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525;
  wire n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557;
  wire n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565;
  wire n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572;
  nand g8 (QUOTIENT[9], n_46, n_49);
  nand g20 (QUOTIENT[7], n_66, n_69);
  nand g32 (QUOTIENT[5], n_94, n_97);
  nand g44 (QUOTIENT[3], n_132, n_135);
  or g55 (QUOTIENT[0], n_186, n_1572);
  xor g57 (n_277, B[0], B[1]);
  nand g58 (n_198, B[0], B[1]);
  nand g63 (n_204, B[1], B[2]);
  nand g9 (n_206, B[2], B[3]);
  nand g11 (n_208, B[3], B[4]);
  nand g65 (n_212, B[4], B[5]);
  nand g67 (n_214, B[5], B[6]);
  nand g69 (n_218, B[6], B[7]);
  nand g71 (n_220, B[7], B[8]);
  nand g21 (n_224, B[8], B[9]);
  nand g74 (n_228, n_204, n_1358);
  nor g75 (n_209, n_206, n_207);
  nor g78 (n_231, n_289, n_207);
  nor g79 (n_215, n_212, n_213);
  nor g34 (n_237, n_291, n_213);
  nor g35 (n_221, n_218, n_219);
  nor g82 (n_239, n_223, n_219);
  nand g45 (n_264, n_206, n_1390);
  nand g46 (n_233, n_231, n_228);
  nand g47 (n_244, n_1362, n_233);
  nor g48 (n_235, n_223, n_234);
  nand g95 (n_252, n_237, n_239);
  nand g98 (n_268, n_212, n_1402);
  nand g99 (n_247, n_237, n_244);
  nand g100 (n_270, n_234, n_247);
  nand g103 (n_273, n_1391, n_1403);
  nand g106 (n_256, n_1392, n_1404);
  nand g109 (n_276, n_224, n_1406);
  nand g110 (n_260, n_1345, n_256);
  xnor g115 (n_32, n_228, n_1359);
  xnor g118 (n_33, n_264, n_1361);
  xnor g120 (n_34, n_244, n_1363);
  xnor g123 (n_35, n_268, n_1364);
  xnor g125 (n_36, n_270, n_1365);
  xnor g128 (n_37, n_273, n_1367);
  xnor g130 (n_38, n_256, n_1369);
  nand g143 (n_286, n_284, n_1375);
  nor g144 (n_289, B[2], B[3]);
  nor g145 (n_291, B[4], B[5]);
  nor g146 (n_223, B[6], B[7]);
  nor g147 (n_307, B[8], B[9]);
  nand g150 (n_290, n_289, n_286);
  nand g153 (n_301, n_291, n_223);
  xnor g165 (n_42, n_282, n_1377);
  nand g191 (n_323, n_321, n_318);
  nor g192 (n_326, B[1], B[2]);
  nor g193 (n_207, B[3], B[4]);
  nor g194 (n_213, B[5], B[6]);
  nor g195 (n_219, B[7], B[8]);
  nand g198 (n_327, n_326, n_323);
  nand g201 (n_340, n_207, n_213);
  nand g245 (n_365, n_363, n_1389);
  nor g246 (n_368, n_31, n_32);
  nor g247 (n_370, n_33, n_34);
  nor g248 (n_372, n_35, n_36);
  nor g249 (n_373, n_37, n_38);
  nor g250 (n_375, n_1408, n_1407);
  nand g253 (n_369, n_368, n_365);
  nand g256 (n_383, n_370, n_372);
  nand g259 (n_393, n_373, n_375);
  xnor g275 (n_43, n_282, n_1393);
  nand g312 (n_420, n_412, n_1379);
  nor g313 (n_417, n_414, n_415);
  nor g316 (n_423, n_419, n_415);
  nand g322 (n_446, n_414, n_1417);
  nand g323 (n_425, n_423, n_420);
  nand g324 (n_429, n_1411, n_425);
  xnor g339 (n_56, n_410, n_1380);
  xnor g341 (n_58, n_420, n_1414);
  xnor g344 (n_61, n_446, n_1418);
  nand g371 (n_469, n_461, n_458);
  nor g372 (n_466, n_463, n_464);
  nor g375 (n_472, n_468, n_464);
  nand g381 (n_499, n_463, n_1419);
  nand g382 (n_474, n_472, n_469);
  nand g383 (n_480, n_1412, n_474);
  xnor g404 (n_59, n_469, n_1415);
  xnor g407 (n_62, n_499, n_1420);
  nand g437 (n_523, n_515, n_1394);
  nor g438 (n_520, n_517, n_518);
  nor g441 (n_526, n_522, n_518);
  nand g448 (n_557, n_517, n_1421);
  nand g449 (n_528, n_526, n_523);
  nand g450 (n_535, n_1413, n_528);
  xnor g472 (n_57, n_410, n_1395);
  xnor g474 (n_60, n_523, n_1416);
  xnor g477 (n_63, n_557, n_1422);
  nand g519 (n_590, n_576, n_1382);
  nor g520 (n_581, n_578, n_579);
  nor g523 (n_593, n_583, n_579);
  nor g524 (n_587, n_584, n_585);
  nor g527 (n_598, n_589, n_585);
  nand g532 (n_620, n_578, n_1436);
  nand g533 (n_595, n_593, n_590);
  nand g534 (n_603, n_1428, n_595);
  nand g540 (n_610, n_598, n_223);
  nand g543 (n_624, n_584, n_1454);
  nand g554 (n_92, n_307, n_1457);
  xnor g556 (n_78, n_574, n_1383);
  xnor g558 (n_80, n_590, n_1433);
  xnor g561 (n_83, n_620, n_1437);
  xnor g563 (n_86, n_603, n_1442);
  xnor g566 (n_89, n_624, n_1445);
  nand g596 (n_656, n_642, n_639);
  nor g597 (n_647, n_644, n_645);
  nor g600 (n_659, n_649, n_645);
  nor g601 (n_653, n_650, n_651);
  nor g604 (n_664, n_655, n_651);
  nand g609 (n_690, n_644, n_1438);
  nand g610 (n_661, n_659, n_656);
  nand g611 (n_671, n_1430, n_661);
  nand g617 (n_678, n_664, n_213);
  nand g622 (n_694, n_650, n_1455);
  xnor g639 (n_81, n_656, n_1434);
  xnor g642 (n_84, n_690, n_1439);
  xnor g644 (n_87, n_671, n_1443);
  xnor g647 (n_90, n_694, n_1446);
  nand g679 (n_727, n_713, n_1396);
  nor g680 (n_718, n_715, n_716);
  nor g683 (n_730, n_720, n_716);
  nor g684 (n_724, n_721, n_722);
  nor g687 (n_735, n_726, n_722);
  nand g693 (n_765, n_715, n_1440);
  nand g694 (n_732, n_730, n_727);
  nand g695 (n_743, n_1432, n_732);
  nand g701 (n_750, n_735, n_372);
  nand g707 (n_769, n_721, n_1456);
  xnor g724 (n_79, n_574, n_1397);
  xnor g726 (n_82, n_727, n_1435);
  xnor g729 (n_85, n_765, n_1441);
  xnor g731 (n_88, n_743, n_1444);
  xnor g734 (n_91, n_769, n_1447);
  nand g780 (n_811, n_791, n_1385);
  nor g781 (n_796, n_793, n_794);
  nor g784 (n_814, n_798, n_794);
  nor g785 (n_802, n_799, n_800);
  nor g788 (n_820, n_804, n_800);
  nor g789 (n_808, n_805, n_806);
  nor g792 (n_822, n_810, n_806);
  nand g796 (n_846, n_793, n_1479);
  nand g797 (n_816, n_814, n_811);
  nand g798 (n_827, n_1462, n_816);
  nor g799 (n_818, n_810, n_817);
  nand g808 (n_835, n_820, n_822);
  nand g811 (n_850, n_799, n_1506);
  nand g812 (n_830, n_820, n_827);
  nand g813 (n_852, n_817, n_830);
  nand g816 (n_855, n_1500, n_1501);
  nand g819 (n_839, n_1494, n_1495);
  nand g822 (n_130, n_307, n_839);
  xnor g824 (n_109, n_789, n_1386);
  xnor g826 (n_112, n_811, n_1476);
  xnor g829 (n_115, n_846, n_1480);
  xnor g831 (n_118, n_827, n_1485);
  xnor g834 (n_121, n_850, n_1488);
  xnor g836 (n_124, n_852, n_1467);
  xnor g839 (n_127, n_855, n_1471);
  nand g871 (n_891, n_871, n_868);
  nor g872 (n_876, n_873, n_874);
  nor g875 (n_894, n_878, n_874);
  nor g876 (n_882, n_879, n_880);
  nor g879 (n_900, n_884, n_880);
  nor g880 (n_888, n_885, n_886);
  nor g883 (n_902, n_890, n_886);
  nand g887 (n_930, n_873, n_1481);
  nand g888 (n_896, n_894, n_891);
  nand g889 (n_909, n_1464, n_896);
  nor g890 (n_898, n_890, n_897);
  nand g899 (n_917, n_900, n_902);
  nand g904 (n_934, n_879, n_1507);
  nand g905 (n_912, n_900, n_909);
  nand g906 (n_936, n_897, n_912);
  nand g909 (n_939, n_1502, n_1503);
  nand g912 (n_921, n_1496, n_1497);
  xnor g921 (n_113, n_891, n_1477);
  xnor g924 (n_116, n_930, n_1482);
  xnor g926 (n_119, n_909, n_1486);
  xnor g929 (n_122, n_934, n_1489);
  xnor g931 (n_125, n_936, n_1468);
  xnor g934 (n_128, n_939, n_1473);
  nand g968 (n_976, n_956, n_1398);
  nor g969 (n_961, n_958, n_959);
  nor g972 (n_979, n_963, n_959);
  nor g973 (n_967, n_964, n_965);
  nor g976 (n_985, n_969, n_965);
  nor g977 (n_973, n_970, n_971);
  nor g980 (n_987, n_975, n_971);
  nand g985 (n_1019, n_958, n_1483);
  nand g986 (n_981, n_979, n_976);
  nand g987 (n_995, n_1466, n_981);
  nor g988 (n_983, n_975, n_982);
  nand g997 (n_1003, n_985, n_987);
  nand g1003 (n_1023, n_964, n_1508);
  nand g1004 (n_998, n_985, n_995);
  nand g1005 (n_1025, n_982, n_998);
  nand g1008 (n_1028, n_1504, n_1505);
  nand g1011 (n_1007, n_1498, n_1499);
  xnor g1020 (n_111, n_789, n_1399);
  xnor g1022 (n_114, n_976, n_1478);
  xnor g1025 (n_117, n_1019, n_1484);
  xnor g1027 (n_120, n_995, n_1487);
  xnor g1030 (n_123, n_1023, n_1490);
  xnor g1032 (n_126, n_1025, n_1469);
  xnor g1035 (n_129, n_1028, n_1475);
  nand g1086 (n_1075, n_1355, n_1388);
  nor g1087 (n_1054, n_1530, n_1052);
  nor g1090 (n_1078, n_1532, n_1052);
  nor g1091 (n_1060, n_1525, n_1058);
  nor g1094 (n_1084, n_1533, n_1058);
  nor g1095 (n_1066, n_1528, n_1064);
  nor g1098 (n_1086, n_1527, n_1064);
  nor g1099 (n_1072, n_1522, n_1070);
  nor g1102 (n_1106, n_1524, n_1070);
  nand g1106 (n_1080, n_1078, n_1075);
  nand g1107 (n_1091, n_1554, n_1080);
  nand g1117 (n_1099, n_1084, n_1086);
  nand g1128 (n_1103, n_1565, n_1566);
  nand g1132 (n_1108, n_1106, n_1103);
  nand g1133 (n_1045, n_1551, n_1108);
  nand g1191 (n_1169, n_1353, n_1354);
  nor g1192 (n_1148, n_1517, n_1146);
  nor g1195 (n_1172, n_1519, n_1146);
  nor g1196 (n_1154, n_1512, n_1152);
  nor g1199 (n_1178, n_1520, n_1152);
  nor g1200 (n_1160, n_1515, n_1158);
  nor g1203 (n_1180, n_1514, n_1158);
  nor g1204 (n_1166, n_1510, n_1164);
  nor g1207 (n_1187, n_1521, n_1164);
  nand g1211 (n_1174, n_1172, n_1169);
  nand g1212 (n_1189, n_1549, n_1174);
  nand g1222 (n_1197, n_1178, n_1180);
  nor g1223 (n_1186, B[9], n_1546);
  nand g1236 (n_1201, n_1563, n_1564);
  nand g1304 (n_1270, n_1373, n_1400);
  nor g1305 (n_1249, n_1541, n_1247);
  nor g1308 (n_1273, n_1543, n_1247);
  nor g1309 (n_1255, n_1536, n_1253);
  nor g1312 (n_1279, n_1544, n_1253);
  nor g1313 (n_1261, n_1539, n_1259);
  nor g1316 (n_1281, n_1538, n_1259);
  nor g1317 (n_1267, n_1534, n_1265);
  nor g1320 (n_1288, n_1545, n_1265);
  nand g1325 (n_1275, n_1273, n_1270);
  nand g1326 (n_1293, n_1558, n_1275);
  nand g1336 (n_1301, n_1279, n_1281);
  nand g1342 (n_1312, n_1288, n_375);
  nand g1353 (n_1305, n_1567, n_1568);
  or g1404 (n_284, B[1], wc);
  not gc (wc, A[9]);
  or g1405 (n_282, wc0, A[8]);
  not gc0 (wc0, B[0]);
  and g1406 (n_1342, B[1], wc1);
  not gc1 (wc1, A[9]);
  or g1407 (n_321, B[0], wc2);
  not gc2 (wc2, A[9]);
  and g1408 (n_318, B[0], wc3);
  not gc3 (wc3, A[9]);
  or g1409 (n_1343, B[9], wc4);
  not gc4 (wc4, n_219);
  and g1410 (n_1344, B[9], wc5);
  not gc5 (wc5, n_224);
  and g1411 (n_1345, B[9], wc6);
  not gc6 (wc6, n_307);
  xnor g1412 (n_1346, A[8], B[0]);
  or g1413 (n_412, B[1], wc7);
  not gc7 (wc7, A[7]);
  or g1414 (n_410, wc8, A[6]);
  not gc8 (wc8, B[0]);
  and g1415 (n_1347, B[1], wc9);
  not gc9 (wc9, A[7]);
  or g1416 (n_461, B[0], wc10);
  not gc10 (wc10, A[7]);
  and g1417 (n_458, B[0], wc11);
  not gc11 (wc11, A[7]);
  xnor g1418 (n_1348, A[6], B[0]);
  or g1419 (n_576, B[1], wc12);
  not gc12 (wc12, A[5]);
  or g1420 (n_574, wc13, A[4]);
  not gc13 (wc13, B[0]);
  and g1421 (n_1349, B[1], wc14);
  not gc14 (wc14, A[5]);
  or g1422 (n_642, B[0], wc15);
  not gc15 (wc15, A[5]);
  and g1423 (n_639, B[0], wc16);
  not gc16 (wc16, A[5]);
  xnor g1424 (n_1350, A[4], B[0]);
  or g1425 (n_791, B[1], wc17);
  not gc17 (wc17, A[3]);
  or g1426 (n_789, wc18, A[2]);
  not gc18 (wc18, B[0]);
  and g1427 (n_1351, B[1], wc19);
  not gc19 (wc19, A[3]);
  or g1428 (n_871, B[0], wc20);
  not gc20 (wc20, A[3]);
  and g1429 (n_868, B[0], wc21);
  not gc21 (wc21, A[3]);
  xnor g1430 (n_1352, A[2], B[0]);
  or g1431 (n_1353, B[0], wc22);
  not gc22 (wc22, A[1]);
  and g1432 (n_1354, B[0], wc23);
  not gc23 (wc23, A[1]);
  or g1433 (n_1355, B[1], wc24);
  not gc24 (wc24, A[1]);
  or g1434 (n_1047, wc25, A[0]);
  not gc25 (wc25, B[0]);
  and g1435 (n_1356, B[1], wc26);
  not gc26 (wc26, A[1]);
  or g1436 (n_1357, n_326, wc27);
  not gc27 (wc27, n_204);
  or g1437 (n_1358, n_198, n_326);
  or g1438 (n_1359, n_289, wc28);
  not gc28 (wc28, n_206);
  or g1439 (n_363, wc29, n_277);
  not gc29 (wc29, A[9]);
  and g1440 (n_1360, wc30, n_277);
  not gc30 (wc30, A[9]);
  or g1441 (n_1361, n_207, wc31);
  not gc31 (wc31, n_208);
  and g1442 (n_1362, wc32, n_208);
  not gc32 (wc32, n_209);
  or g1443 (n_1363, n_291, wc33);
  not gc33 (wc33, n_212);
  or g1444 (n_1364, n_213, wc34);
  not gc34 (wc34, n_214);
  and g1445 (n_234, wc35, n_214);
  not gc35 (wc35, n_215);
  or g1446 (n_1365, n_223, wc36);
  not gc36 (wc36, n_218);
  or g1447 (n_1366, n_223, wc37);
  not gc37 (wc37, n_237);
  or g1448 (n_1367, n_219, wc38);
  not gc38 (wc38, n_220);
  and g1449 (n_1368, wc39, n_220);
  not gc39 (wc39, n_221);
  or g1450 (n_1369, n_307, wc40);
  not gc40 (wc40, n_224);
  or g1451 (n_515, wc41, n_277);
  not gc41 (wc41, A[7]);
  and g1452 (n_1370, wc42, n_277);
  not gc42 (wc42, A[7]);
  or g1453 (n_713, wc43, n_277);
  not gc43 (wc43, A[5]);
  and g1454 (n_1371, wc44, n_277);
  not gc44 (wc44, A[5]);
  or g1455 (n_956, wc45, n_277);
  not gc45 (wc45, A[3]);
  and g1456 (n_1372, wc46, n_277);
  not gc46 (wc46, A[3]);
  or g1457 (n_1373, wc47, n_277);
  not gc47 (wc47, A[1]);
  and g1458 (n_1374, wc48, n_277);
  not gc48 (wc48, A[1]);
  or g1459 (n_1375, n_1342, wc49);
  not gc49 (wc49, n_282);
  xor g1460 (n_31, n_198, n_1357);
  and g1461 (n_1376, wc50, n_239);
  not gc50 (wc50, n_234);
  or g1462 (n_1377, n_1342, wc51);
  not gc51 (wc51, n_284);
  or g1463 (n_1378, n_318, wc52);
  not gc52 (wc52, n_321);
  or g1464 (n_1379, n_1347, wc53);
  not gc53 (wc53, n_410);
  or g1465 (n_1380, n_1347, wc54);
  not gc54 (wc54, n_412);
  or g1466 (n_1381, n_458, wc55);
  not gc55 (wc55, n_461);
  or g1467 (n_1382, n_1349, wc56);
  not gc56 (wc56, n_574);
  or g1468 (n_1383, n_1349, wc57);
  not gc57 (wc57, n_576);
  or g1469 (n_1384, n_639, wc58);
  not gc58 (wc58, n_642);
  or g1470 (n_1385, n_1351, wc59);
  not gc59 (wc59, n_789);
  or g1471 (n_1386, n_1351, wc60);
  not gc60 (wc60, n_791);
  or g1472 (n_1387, n_868, wc61);
  not gc61 (wc61, n_871);
  or g1473 (n_1388, n_1356, wc62);
  not gc62 (wc62, n_1047);
  or g1474 (n_1389, n_1360, wc63);
  not gc63 (wc63, n_282);
  or g1475 (n_1390, n_289, wc64);
  not gc64 (wc64, n_228);
  and g1476 (n_1391, wc65, n_218);
  not gc65 (wc65, n_235);
  and g1477 (n_1392, wc66, n_1368);
  not gc66 (wc66, n_1376);
  or g1478 (n_1393, n_1360, wc67);
  not gc67 (wc67, n_363);
  or g1479 (n_1394, n_1370, wc68);
  not gc68 (wc68, n_410);
  or g1480 (n_1395, n_1370, wc69);
  not gc69 (wc69, n_515);
  or g1481 (n_1396, n_1371, wc70);
  not gc70 (wc70, n_574);
  or g1482 (n_1397, n_1371, wc71);
  not gc71 (wc71, n_713);
  or g1483 (n_1398, n_1372, wc72);
  not gc72 (wc72, n_789);
  or g1484 (n_1399, n_1372, wc73);
  not gc73 (wc73, n_956);
  or g1485 (n_1400, n_1374, wc74);
  not gc74 (wc74, n_1047);
  or g1486 (n_1401, n_327, n_340);
  or g1487 (n_1402, n_291, wc75);
  not gc75 (wc75, n_244);
  or g1488 (n_1403, n_1366, wc76);
  not gc76 (wc76, n_244);
  or g1489 (n_1404, n_252, wc77);
  not gc77 (wc77, n_244);
  or g1490 (n_1405, n_290, n_301);
  or g1491 (n_46, n_1343, n_1401);
  or g1492 (n_1406, n_307, wc78);
  not gc78 (wc78, n_256);
  or g1493 (n_44, n_1405, wc79);
  not gc79 (wc79, n_307);
  or g1494 (n_1407, n_1344, wc80);
  not gc80 (wc80, n_260);
  xor g1495 (n_1408, n_276, B[9]);
  and g1496 (n_47, wc81, n_46);
  not gc81 (wc81, n_44);
  or g1497 (n_1409, n_369, n_383);
  or g1498 (n_49, n_393, n_1409);
  and g1499 (n_50, n_49, wc82);
  not gc82 (wc82, n_46);
  or g1500 (QUOTIENT[8], wc83, n_47);
  not gc83 (wc83, n_49);
  or g1501 (n_53, wc84, wc85, wc87, wc88);
  and gc90 (wc88, wc89, wc90);
  not gc89 (wc90, n_1346);
  not gc88 (wc89, n_49);
  and gc87 (wc87, A[8], n_50);
  and gc86 (wc85, n_47, wc86);
  not gc85 (wc86, n_1346);
  and gc84 (wc84, A[8], n_44);
  or g1502 (n_54, wc91, wc92, wc93, wc94);
  and gc95 (wc94, wc95, n_43);
  not gc94 (wc95, n_49);
  and gc93 (wc93, n_50, n_1378);
  and gc92 (wc92, n_47, n_42);
  and gc91 (wc91, A[9], n_44);
  or g1503 (n_414, B[2], wc96);
  not gc96 (wc96, n_53);
  and g1504 (n_415, B[3], wc97);
  not gc97 (wc97, n_54);
  or g1505 (n_416, B[3], wc98);
  not gc98 (wc98, n_54);
  and g1506 (n_419, B[2], wc99);
  not gc99 (wc99, n_53);
  or g1507 (n_463, B[1], wc100);
  not gc100 (wc100, n_53);
  and g1508 (n_464, B[2], wc101);
  not gc101 (wc101, n_54);
  or g1509 (n_465, B[2], wc102);
  not gc102 (wc102, n_54);
  and g1510 (n_468, B[1], wc103);
  not gc103 (wc103, n_53);
  or g1511 (n_517, wc104, n_31);
  not gc104 (wc104, n_53);
  and g1512 (n_518, wc105, n_32);
  not gc105 (wc105, n_54);
  or g1513 (n_519, wc106, n_32);
  not gc106 (wc106, n_54);
  and g1514 (n_522, wc107, n_31);
  not gc107 (wc107, n_53);
  and g1515 (n_1411, n_416, wc108);
  not gc108 (wc108, n_417);
  and g1516 (n_1412, n_465, wc109);
  not gc109 (wc109, n_466);
  and g1517 (n_1413, n_519, wc110);
  not gc110 (wc110, n_520);
  or g1518 (n_1414, n_419, wc111);
  not gc111 (wc111, n_414);
  or g1519 (n_1415, n_468, wc112);
  not gc112 (wc112, n_463);
  or g1520 (n_1416, n_522, wc113);
  not gc113 (wc113, n_517);
  or g1521 (n_1417, n_419, wc114);
  not gc114 (wc114, n_420);
  or g1522 (n_1418, wc115, n_415);
  not gc115 (wc115, n_416);
  or g1523 (n_1419, n_468, wc116);
  not gc116 (wc116, n_469);
  or g1524 (n_1420, wc117, n_464);
  not gc117 (wc117, n_465);
  or g1525 (n_1421, n_522, wc118);
  not gc118 (wc118, n_523);
  or g1526 (n_1422, wc119, n_518);
  not gc119 (wc119, n_519);
  or g1527 (n_1423, wc120, n_301);
  not gc120 (wc120, n_429);
  or g1528 (n_1424, wc121, n_340);
  not gc121 (wc121, n_480);
  or g1529 (n_1425, wc122, n_383);
  not gc122 (wc122, n_535);
  or g1530 (n_64, n_1423, wc123);
  not gc123 (wc123, n_307);
  or g1531 (n_66, n_1343, n_1424);
  or g1532 (n_69, n_393, n_1425);
  and g1533 (n_67, n_66, wc124);
  not gc124 (wc124, n_64);
  and g1534 (n_70, n_69, wc125);
  not gc125 (wc125, n_66);
  or g1535 (QUOTIENT[6], n_67, wc126);
  not gc126 (wc126, n_69);
  or g1536 (n_75, wc127, wc128, wc129, wc130);
  and gc131 (wc130, wc131, n_60);
  not gc130 (wc131, n_69);
  and gc129 (wc129, n_70, n_59);
  and gc128 (wc128, n_67, n_58);
  and gc127 (wc127, n_64, n_53);
  or g1537 (n_76, wc132, wc133, wc134, wc135);
  and gc136 (wc135, wc136, n_63);
  not gc135 (wc136, n_69);
  and gc134 (wc134, n_70, n_62);
  and gc133 (wc133, n_67, n_61);
  and gc132 (wc132, n_64, n_54);
  or g1538 (n_73, wc137, wc138, wc140, wc141);
  and gc143 (wc141, wc142, wc143);
  not gc142 (wc143, n_1348);
  not gc141 (wc142, n_69);
  and gc140 (wc140, A[6], n_70);
  and gc139 (wc138, n_67, wc139);
  not gc138 (wc139, n_1348);
  and gc137 (wc137, A[6], n_64);
  or g1539 (n_74, wc144, wc145, wc146, wc147);
  and gc148 (wc147, wc148, n_57);
  not gc147 (wc148, n_69);
  and gc146 (wc146, n_70, n_1381);
  and gc145 (wc145, n_67, n_56);
  and gc144 (wc144, A[7], n_64);
  or g1540 (n_584, B[4], wc149);
  not gc149 (wc149, n_75);
  and g1541 (n_585, B[5], wc150);
  not gc150 (wc150, n_76);
  or g1542 (n_586, B[5], wc151);
  not gc151 (wc151, n_76);
  or g1543 (n_578, B[2], wc152);
  not gc152 (wc152, n_73);
  and g1544 (n_579, B[3], wc153);
  not gc153 (wc153, n_74);
  or g1545 (n_580, B[3], wc154);
  not gc154 (wc154, n_74);
  and g1546 (n_583, B[2], wc155);
  not gc155 (wc155, n_73);
  and g1547 (n_589, B[4], wc156);
  not gc156 (wc156, n_75);
  or g1548 (n_650, B[3], wc157);
  not gc157 (wc157, n_75);
  and g1549 (n_651, B[4], wc158);
  not gc158 (wc158, n_76);
  or g1550 (n_652, B[4], wc159);
  not gc159 (wc159, n_76);
  or g1551 (n_644, B[1], wc160);
  not gc160 (wc160, n_73);
  and g1552 (n_645, B[2], wc161);
  not gc161 (wc161, n_74);
  or g1553 (n_646, B[2], wc162);
  not gc162 (wc162, n_74);
  and g1554 (n_649, B[1], wc163);
  not gc163 (wc163, n_73);
  and g1555 (n_655, B[3], wc164);
  not gc164 (wc164, n_75);
  or g1556 (n_721, wc165, n_33);
  not gc165 (wc165, n_75);
  and g1557 (n_722, wc166, n_34);
  not gc166 (wc166, n_76);
  or g1558 (n_723, wc167, n_34);
  not gc167 (wc167, n_76);
  or g1559 (n_715, wc168, n_31);
  not gc168 (wc168, n_73);
  and g1560 (n_716, wc169, n_32);
  not gc169 (wc169, n_74);
  or g1561 (n_717, wc170, n_32);
  not gc170 (wc170, n_74);
  and g1562 (n_720, wc171, n_31);
  not gc171 (wc171, n_73);
  and g1563 (n_726, wc172, n_33);
  not gc172 (wc172, n_75);
  and g1564 (n_1427, n_586, wc173);
  not gc173 (wc173, n_587);
  and g1565 (n_1428, n_580, wc174);
  not gc174 (wc174, n_581);
  and g1566 (n_1429, n_652, wc175);
  not gc175 (wc175, n_653);
  and g1567 (n_1430, n_646, wc176);
  not gc176 (wc176, n_647);
  and g1568 (n_1431, n_723, wc177);
  not gc177 (wc177, n_724);
  and g1569 (n_1432, n_717, wc178);
  not gc178 (wc178, n_718);
  or g1570 (n_1433, n_583, wc179);
  not gc179 (wc179, n_578);
  or g1571 (n_1434, n_649, wc180);
  not gc180 (wc180, n_644);
  or g1572 (n_1435, n_720, wc181);
  not gc181 (wc181, n_715);
  or g1573 (n_1436, n_583, wc182);
  not gc182 (wc182, n_590);
  or g1574 (n_1437, wc183, n_579);
  not gc183 (wc183, n_580);
  or g1575 (n_1438, n_649, wc184);
  not gc184 (wc184, n_656);
  or g1576 (n_1439, wc185, n_645);
  not gc185 (wc185, n_646);
  or g1577 (n_1440, n_720, wc186);
  not gc186 (wc186, n_727);
  or g1578 (n_1441, wc187, n_716);
  not gc187 (wc187, n_717);
  or g1579 (n_1442, n_589, wc188);
  not gc188 (wc188, n_584);
  or g1580 (n_1443, n_655, wc189);
  not gc189 (wc189, n_650);
  or g1581 (n_1444, n_726, wc190);
  not gc190 (wc190, n_721);
  or g1582 (n_1445, wc191, n_585);
  not gc191 (wc191, n_586);
  or g1583 (n_1446, wc192, n_651);
  not gc192 (wc192, n_652);
  or g1584 (n_1447, wc193, n_722);
  not gc193 (wc193, n_723);
  and g1585 (n_1448, wc194, n_223);
  not gc194 (wc194, n_1427);
  and g1586 (n_1449, wc195, n_213);
  not gc195 (wc195, n_1429);
  and g1587 (n_1450, wc196, n_372);
  not gc196 (wc196, n_1431);
  or g1588 (n_1451, n_610, wc197);
  not gc197 (wc197, n_603);
  or g1589 (n_1452, n_678, wc198);
  not gc198 (wc198, n_671);
  or g1590 (n_1453, n_750, wc199);
  not gc199 (wc199, n_743);
  or g1591 (n_1454, n_589, wc200);
  not gc200 (wc200, n_603);
  or g1592 (n_1455, n_655, wc201);
  not gc201 (wc201, n_671);
  or g1593 (n_1456, n_726, wc202);
  not gc202 (wc202, n_743);
  or g1594 (n_1457, wc203, n_1448);
  not gc203 (wc203, n_1451);
  or g1595 (n_1458, wc204, n_1449);
  not gc204 (wc204, n_1452);
  or g1596 (n_1459, wc205, n_1450);
  not gc205 (wc205, n_1453);
  or g1597 (n_94, wc206, n_1343);
  not gc206 (wc206, n_1458);
  or g1598 (n_97, wc207, n_393);
  not gc207 (wc207, n_1459);
  and g1599 (n_95, n_94, wc208);
  not gc208 (wc208, n_92);
  and g1600 (n_98, n_97, wc209);
  not gc209 (wc209, n_94);
  or g1601 (QUOTIENT[4], n_95, wc210);
  not gc210 (wc210, n_97);
  or g1602 (n_103, wc211, wc212, wc213, wc214);
  and gc215 (wc214, wc215, n_82);
  not gc214 (wc215, n_97);
  and gc213 (wc213, n_98, n_81);
  and gc212 (wc212, n_95, n_80);
  and gc211 (wc211, n_73, n_92);
  or g1603 (n_104, wc216, wc217, wc218, wc219);
  and gc220 (wc219, wc220, n_85);
  not gc219 (wc220, n_97);
  and gc218 (wc218, n_98, n_84);
  and gc217 (wc217, n_95, n_83);
  and gc216 (wc216, n_74, n_92);
  or g1604 (n_105, wc221, wc222, wc223, wc224);
  and gc225 (wc224, wc225, n_88);
  not gc224 (wc225, n_97);
  and gc223 (wc223, n_98, n_87);
  and gc222 (wc222, n_95, n_86);
  and gc221 (wc221, n_75, n_92);
  or g1605 (n_106, wc226, wc227, wc228, wc229);
  and gc230 (wc229, wc230, n_91);
  not gc229 (wc230, n_97);
  and gc228 (wc228, n_98, n_90);
  and gc227 (wc227, n_95, n_89);
  and gc226 (wc226, n_76, n_92);
  or g1606 (n_101, wc231, wc232, wc234, wc235);
  and gc237 (wc235, wc236, wc237);
  not gc236 (wc237, n_1350);
  not gc235 (wc236, n_97);
  and gc234 (wc234, A[4], n_98);
  and gc233 (wc232, n_95, wc233);
  not gc232 (wc233, n_1350);
  and gc231 (wc231, A[4], n_92);
  or g1607 (n_102, wc238, wc239, wc240, wc241);
  and gc242 (wc241, wc242, n_79);
  not gc241 (wc242, n_97);
  and gc240 (wc240, n_98, n_1384);
  and gc239 (wc239, n_95, n_78);
  and gc238 (wc238, A[5], n_92);
  or g1608 (n_799, B[4], wc243);
  not gc243 (wc243, n_103);
  and g1609 (n_800, B[5], wc244);
  not gc244 (wc244, n_104);
  or g1610 (n_801, B[5], wc245);
  not gc245 (wc245, n_104);
  and g1611 (n_810, B[6], wc246);
  not gc246 (wc246, n_105);
  and g1612 (n_806, B[7], wc247);
  not gc247 (wc247, n_106);
  or g1613 (n_805, B[6], wc248);
  not gc248 (wc248, n_105);
  or g1614 (n_807, B[7], wc249);
  not gc249 (wc249, n_106);
  or g1615 (n_793, B[2], wc250);
  not gc250 (wc250, n_101);
  and g1616 (n_794, B[3], wc251);
  not gc251 (wc251, n_102);
  or g1617 (n_795, B[3], wc252);
  not gc252 (wc252, n_102);
  and g1618 (n_798, B[2], wc253);
  not gc253 (wc253, n_101);
  and g1619 (n_804, B[4], wc254);
  not gc254 (wc254, n_103);
  or g1620 (n_879, B[3], wc255);
  not gc255 (wc255, n_103);
  and g1621 (n_880, B[4], wc256);
  not gc256 (wc256, n_104);
  or g1622 (n_881, B[4], wc257);
  not gc257 (wc257, n_104);
  and g1623 (n_890, B[5], wc258);
  not gc258 (wc258, n_105);
  and g1624 (n_886, B[6], wc259);
  not gc259 (wc259, n_106);
  or g1625 (n_885, B[5], wc260);
  not gc260 (wc260, n_105);
  or g1626 (n_887, B[6], wc261);
  not gc261 (wc261, n_106);
  or g1627 (n_873, B[1], wc262);
  not gc262 (wc262, n_101);
  and g1628 (n_874, B[2], wc263);
  not gc263 (wc263, n_102);
  or g1629 (n_875, B[2], wc264);
  not gc264 (wc264, n_102);
  and g1630 (n_878, B[1], wc265);
  not gc265 (wc265, n_101);
  and g1631 (n_884, B[3], wc266);
  not gc266 (wc266, n_103);
  or g1632 (n_964, wc267, n_33);
  not gc267 (wc267, n_103);
  and g1633 (n_965, wc268, n_34);
  not gc268 (wc268, n_104);
  or g1634 (n_966, wc269, n_34);
  not gc269 (wc269, n_104);
  and g1635 (n_975, wc270, n_35);
  not gc270 (wc270, n_105);
  and g1636 (n_971, wc271, n_36);
  not gc271 (wc271, n_106);
  or g1637 (n_970, wc272, n_35);
  not gc272 (wc272, n_105);
  or g1638 (n_972, wc273, n_36);
  not gc273 (wc273, n_106);
  or g1639 (n_958, wc274, n_31);
  not gc274 (wc274, n_101);
  and g1640 (n_959, wc275, n_32);
  not gc275 (wc275, n_102);
  or g1641 (n_960, wc276, n_32);
  not gc276 (wc276, n_102);
  and g1642 (n_963, wc277, n_31);
  not gc277 (wc277, n_101);
  and g1643 (n_969, wc278, n_33);
  not gc278 (wc278, n_103);
  and g1644 (n_817, n_801, wc279);
  not gc279 (wc279, n_802);
  and g1645 (n_1461, n_807, wc280);
  not gc280 (wc280, n_808);
  and g1646 (n_1462, n_795, wc281);
  not gc281 (wc281, n_796);
  and g1647 (n_897, n_881, wc282);
  not gc282 (wc282, n_882);
  and g1648 (n_1463, n_887, wc283);
  not gc283 (wc283, n_888);
  and g1649 (n_1464, n_875, wc284);
  not gc284 (wc284, n_876);
  and g1650 (n_982, n_966, wc285);
  not gc285 (wc285, n_967);
  and g1651 (n_1465, n_972, wc286);
  not gc286 (wc286, n_973);
  and g1652 (n_1466, n_960, wc287);
  not gc287 (wc287, n_961);
  or g1653 (n_1467, wc288, n_810);
  not gc288 (wc288, n_805);
  or g1654 (n_1468, wc289, n_890);
  not gc289 (wc289, n_885);
  or g1655 (n_1469, wc290, n_975);
  not gc290 (wc290, n_970);
  or g1656 (n_1470, n_810, wc291);
  not gc291 (wc291, n_820);
  or g1657 (n_1471, wc292, n_806);
  not gc292 (wc292, n_807);
  or g1658 (n_1472, n_890, wc293);
  not gc293 (wc293, n_900);
  or g1659 (n_1473, wc294, n_886);
  not gc294 (wc294, n_887);
  or g1660 (n_1474, n_975, wc295);
  not gc295 (wc295, n_985);
  or g1661 (n_1475, wc296, n_971);
  not gc296 (wc296, n_972);
  or g1662 (n_1476, n_798, wc297);
  not gc297 (wc297, n_793);
  or g1663 (n_1477, n_878, wc298);
  not gc298 (wc298, n_873);
  or g1664 (n_1478, n_963, wc299);
  not gc299 (wc299, n_958);
  or g1665 (n_1479, n_798, wc300);
  not gc300 (wc300, n_811);
  or g1666 (n_1480, wc301, n_794);
  not gc301 (wc301, n_795);
  or g1667 (n_1481, n_878, wc302);
  not gc302 (wc302, n_891);
  or g1668 (n_1482, wc303, n_874);
  not gc303 (wc303, n_875);
  or g1669 (n_1483, n_963, wc304);
  not gc304 (wc304, n_976);
  or g1670 (n_1484, wc305, n_959);
  not gc305 (wc305, n_960);
  or g1671 (n_1485, n_804, wc306);
  not gc306 (wc306, n_799);
  or g1672 (n_1486, n_884, wc307);
  not gc307 (wc307, n_879);
  or g1673 (n_1487, n_969, wc308);
  not gc308 (wc308, n_964);
  or g1674 (n_1488, wc309, n_800);
  not gc309 (wc309, n_801);
  or g1675 (n_1489, wc310, n_880);
  not gc310 (wc310, n_881);
  or g1676 (n_1490, wc311, n_965);
  not gc311 (wc311, n_966);
  and g1677 (n_1491, wc312, n_822);
  not gc312 (wc312, n_817);
  and g1678 (n_1492, wc313, n_902);
  not gc313 (wc313, n_897);
  and g1679 (n_1493, wc314, n_987);
  not gc314 (wc314, n_982);
  and g1680 (n_1494, wc315, n_1461);
  not gc315 (wc315, n_1491);
  or g1681 (n_1495, n_835, wc316);
  not gc316 (wc316, n_827);
  and g1682 (n_1496, wc317, n_1463);
  not gc317 (wc317, n_1492);
  or g1683 (n_1497, n_917, wc318);
  not gc318 (wc318, n_909);
  and g1684 (n_1498, wc319, n_1465);
  not gc319 (wc319, n_1493);
  or g1685 (n_1499, n_1003, wc320);
  not gc320 (wc320, n_995);
  and g1686 (n_1500, n_805, wc321);
  not gc321 (wc321, n_818);
  or g1687 (n_1501, n_1470, wc322);
  not gc322 (wc322, n_827);
  and g1688 (n_1502, n_885, wc323);
  not gc323 (wc323, n_898);
  or g1689 (n_1503, n_1472, wc324);
  not gc324 (wc324, n_909);
  and g1690 (n_1504, n_970, wc325);
  not gc325 (wc325, n_983);
  or g1691 (n_1505, n_1474, wc326);
  not gc326 (wc326, n_995);
  or g1692 (n_1506, n_804, wc327);
  not gc327 (wc327, n_827);
  or g1693 (n_1507, n_884, wc328);
  not gc328 (wc328, n_909);
  or g1694 (n_1508, n_969, wc329);
  not gc329 (wc329, n_995);
  or g1695 (n_132, n_1343, wc330);
  not gc330 (wc330, n_921);
  or g1696 (n_135, wc331, n_393);
  not gc331 (wc331, n_1007);
  and g1697 (n_133, n_132, wc332);
  not gc332 (wc332, n_130);
  and g1698 (n_136, n_135, wc333);
  not gc333 (wc333, n_132);
  or g1699 (QUOTIENT[2], n_133, wc334);
  not gc334 (wc334, n_135);
  or g1700 (n_147, wc335, wc336, wc337, wc338);
  and gc339 (wc338, wc339, n_126);
  not gc338 (wc339, n_135);
  and gc337 (wc337, n_136, n_125);
  and gc336 (wc336, n_133, n_124);
  and gc335 (wc335, n_105, n_130);
  or g1701 (n_148, wc340, wc341, wc342, wc343);
  and gc344 (wc343, wc344, n_129);
  not gc343 (wc344, n_135);
  and gc342 (wc342, n_136, n_128);
  and gc341 (wc341, n_133, n_127);
  and gc340 (wc340, n_106, n_130);
  or g1702 (n_143, wc345, wc346, wc347, wc348);
  and gc349 (wc348, wc349, n_114);
  not gc348 (wc349, n_135);
  and gc347 (wc347, n_136, n_113);
  and gc346 (wc346, n_133, n_112);
  and gc345 (wc345, n_101, n_130);
  or g1703 (n_144, wc350, wc351, wc352, wc353);
  and gc354 (wc353, wc354, n_117);
  not gc353 (wc354, n_135);
  and gc352 (wc352, n_136, n_116);
  and gc351 (wc351, n_133, n_115);
  and gc350 (wc350, n_102, n_130);
  or g1704 (n_145, wc355, wc356, wc357, wc358);
  and gc359 (wc358, wc359, n_120);
  not gc358 (wc359, n_135);
  and gc357 (wc357, n_136, n_119);
  and gc356 (wc356, n_133, n_118);
  and gc355 (wc355, n_103, n_130);
  or g1705 (n_146, wc360, wc361, wc362, wc363);
  and gc364 (wc363, wc364, n_123);
  not gc363 (wc364, n_135);
  and gc362 (wc362, n_136, n_122);
  and gc361 (wc361, n_133, n_121);
  and gc360 (wc360, n_104, n_130);
  or g1706 (n_141, wc365, wc366, wc368, wc369);
  and gc371 (wc369, wc370, wc371);
  not gc370 (wc371, n_1352);
  not gc369 (wc370, n_135);
  and gc368 (wc368, A[2], n_136);
  and gc367 (wc366, n_133, wc367);
  not gc366 (wc367, n_1352);
  and gc365 (wc365, A[2], n_130);
  or g1707 (n_142, wc372, wc373, wc374, wc375);
  and gc376 (wc375, wc376, n_111);
  not gc375 (wc376, n_135);
  and gc374 (wc374, n_136, n_1387);
  and gc373 (wc373, n_133, n_109);
  and gc372 (wc372, A[3], n_130);
  or g1708 (n_1510, B[7], wc377);
  not gc377 (wc377, n_147);
  and g1709 (n_1164, B[8], wc378);
  not gc378 (wc378, n_148);
  or g1710 (n_1511, B[8], wc379);
  not gc379 (wc379, n_148);
  or g1711 (n_1512, B[3], wc380);
  not gc380 (wc380, n_143);
  and g1712 (n_1152, B[4], wc381);
  not gc381 (wc381, n_144);
  or g1713 (n_1513, B[4], wc382);
  not gc382 (wc382, n_144);
  and g1714 (n_1514, B[5], wc383);
  not gc383 (wc383, n_145);
  and g1715 (n_1158, B[6], wc384);
  not gc384 (wc384, n_146);
  or g1716 (n_1515, B[5], wc385);
  not gc385 (wc385, n_145);
  or g1717 (n_1516, B[6], wc386);
  not gc386 (wc386, n_146);
  or g1718 (n_1517, B[1], wc387);
  not gc387 (wc387, n_141);
  and g1719 (n_1146, B[2], wc388);
  not gc388 (wc388, n_142);
  or g1720 (n_1518, B[2], wc389);
  not gc389 (wc389, n_142);
  and g1721 (n_1519, B[1], wc390);
  not gc390 (wc390, n_141);
  and g1722 (n_1520, B[3], wc391);
  not gc391 (wc391, n_143);
  and g1723 (n_1521, B[7], wc392);
  not gc392 (wc392, n_147);
  or g1724 (n_1522, B[8], wc393);
  not gc393 (wc393, n_147);
  and g1725 (n_1070, B[9], wc394);
  not gc394 (wc394, n_148);
  or g1726 (n_1523, B[9], wc395);
  not gc395 (wc395, n_148);
  and g1727 (n_1524, B[8], wc396);
  not gc396 (wc396, n_147);
  or g1728 (n_1525, B[4], wc397);
  not gc397 (wc397, n_143);
  and g1729 (n_1058, B[5], wc398);
  not gc398 (wc398, n_144);
  or g1730 (n_1526, B[5], wc399);
  not gc399 (wc399, n_144);
  and g1731 (n_1527, B[6], wc400);
  not gc400 (wc400, n_145);
  and g1732 (n_1064, B[7], wc401);
  not gc401 (wc401, n_146);
  or g1733 (n_1528, B[6], wc402);
  not gc402 (wc402, n_145);
  or g1734 (n_1529, B[7], wc403);
  not gc403 (wc403, n_146);
  or g1735 (n_1530, B[2], wc404);
  not gc404 (wc404, n_141);
  and g1736 (n_1052, B[3], wc405);
  not gc405 (wc405, n_142);
  or g1737 (n_1531, B[3], wc406);
  not gc406 (wc406, n_142);
  and g1738 (n_1532, B[2], wc407);
  not gc407 (wc407, n_141);
  and g1739 (n_1533, B[4], wc408);
  not gc408 (wc408, n_143);
  or g1740 (n_1534, wc409, n_37);
  not gc409 (wc409, n_147);
  and g1741 (n_1265, wc410, n_38);
  not gc410 (wc410, n_148);
  or g1742 (n_1535, wc411, n_38);
  not gc411 (wc411, n_148);
  or g1743 (n_1536, wc412, n_33);
  not gc412 (wc412, n_143);
  and g1744 (n_1253, wc413, n_34);
  not gc413 (wc413, n_144);
  or g1745 (n_1537, wc414, n_34);
  not gc414 (wc414, n_144);
  and g1746 (n_1538, wc415, n_35);
  not gc415 (wc415, n_145);
  and g1747 (n_1259, wc416, n_36);
  not gc416 (wc416, n_146);
  or g1748 (n_1539, wc417, n_35);
  not gc417 (wc417, n_145);
  or g1749 (n_1540, wc418, n_36);
  not gc418 (wc418, n_146);
  or g1750 (n_1541, wc419, n_31);
  not gc419 (wc419, n_141);
  and g1751 (n_1247, wc420, n_32);
  not gc420 (wc420, n_142);
  or g1752 (n_1542, wc421, n_32);
  not gc421 (wc421, n_142);
  and g1753 (n_1543, wc422, n_31);
  not gc422 (wc422, n_141);
  and g1754 (n_1544, wc423, n_33);
  not gc423 (wc423, n_143);
  and g1755 (n_1545, wc424, n_37);
  not gc424 (wc424, n_147);
  and g1756 (n_1546, n_1511, wc425);
  not gc425 (wc425, n_1166);
  and g1757 (n_1547, n_1513, wc426);
  not gc426 (wc426, n_1154);
  and g1758 (n_1548, n_1516, wc427);
  not gc427 (wc427, n_1160);
  and g1759 (n_1549, n_1518, wc428);
  not gc428 (wc428, n_1148);
  or g1760 (n_1550, B[9], wc429);
  not gc429 (wc429, n_1187);
  and g1761 (n_1551, n_1523, wc430);
  not gc430 (wc430, n_1072);
  and g1762 (n_1552, n_1526, wc431);
  not gc431 (wc431, n_1060);
  and g1763 (n_1553, n_1529, wc432);
  not gc432 (wc432, n_1066);
  and g1764 (n_1554, n_1531, wc433);
  not gc433 (wc433, n_1054);
  and g1765 (n_1555, n_1535, wc434);
  not gc434 (wc434, n_1267);
  and g1766 (n_1556, n_1537, wc435);
  not gc435 (wc435, n_1255);
  and g1767 (n_1557, n_1540, wc436);
  not gc436 (wc436, n_1261);
  and g1768 (n_1558, n_1542, wc437);
  not gc437 (wc437, n_1249);
  and g1769 (n_1559, wc438, n_1180);
  not gc438 (wc438, n_1547);
  and g1770 (n_1560, wc439, n_1086);
  not gc439 (wc439, n_1552);
  and g1771 (n_1561, wc440, n_375);
  not gc440 (wc440, n_1555);
  and g1772 (n_1562, wc441, n_1281);
  not gc441 (wc441, n_1556);
  and g1773 (n_1563, wc442, n_1548);
  not gc442 (wc442, n_1559);
  or g1774 (n_1564, n_1197, wc443);
  not gc443 (wc443, n_1189);
  and g1775 (n_1565, wc444, n_1553);
  not gc444 (wc444, n_1560);
  or g1776 (n_1566, n_1099, wc445);
  not gc445 (wc445, n_1091);
  and g1777 (n_1567, wc446, n_1557);
  not gc446 (wc446, n_1562);
  or g1778 (n_1568, n_1301, wc447);
  not gc447 (wc447, n_1293);
  or g1779 (n_1569, n_1550, wc448);
  not gc448 (wc448, n_1201);
  or g1780 (n_1570, wc449, n_1312);
  not gc449 (wc449, n_1305);
  or g1781 (n_1571, wc450, n_1186);
  not gc450 (wc450, n_1569);
  or g1782 (n_186, wc451, n_1561);
  not gc451 (wc451, n_1570);
  and g1783 (n_1572, wc452, n_1045);
  not gc452 (wc452, n_1571);
  or g1784 (QUOTIENT[1], n_1571, n_186);
endmodule

module divide_unsigned_GENERIC(A, B, QUOTIENT);
  input [9:0] A, B;
  output [9:0] QUOTIENT;
  wire [9:0] A, B;
  wire [9:0] QUOTIENT;
  divide_unsigned_GENERIC_REAL g1(.A (A), .B (B), .QUOTIENT (QUOTIENT));
endmodule

module divide_unsigned_16_GENERIC_REAL(A, B, QUOTIENT);
// synthesis_equation "assign QUOTIENT = A / B;"
  input [9:0] A, B;
  output [9:0] QUOTIENT;
  wire [9:0] A, B;
  wire [9:0] QUOTIENT;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_42, n_43, n_44, n_46, n_47, n_49, n_50, n_53;
  wire n_54, n_56, n_57, n_58, n_59, n_60, n_61, n_62;
  wire n_63, n_64, n_66, n_67, n_69, n_70, n_73, n_74;
  wire n_75, n_76, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_94, n_95, n_97, n_98, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_109, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_132, n_133, n_135, n_136, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_186, n_198, n_204, n_206;
  wire n_207, n_208, n_209, n_212, n_213, n_214, n_215, n_218;
  wire n_219, n_220, n_221, n_223, n_224, n_228, n_231, n_233;
  wire n_234, n_235, n_237, n_239, n_244, n_247, n_252, n_256;
  wire n_260, n_264, n_268, n_270, n_273, n_276, n_277, n_282;
  wire n_284, n_286, n_289, n_290, n_291, n_301, n_307, n_318;
  wire n_321, n_323, n_326, n_327, n_340, n_363, n_365, n_368;
  wire n_369, n_370, n_372, n_373, n_375, n_383, n_393, n_410;
  wire n_412, n_414, n_415, n_416, n_417, n_419, n_420, n_423;
  wire n_425, n_429, n_446, n_458, n_461, n_463, n_464, n_465;
  wire n_466, n_468, n_469, n_472, n_474, n_480, n_499, n_515;
  wire n_517, n_518, n_519, n_520, n_522, n_523, n_526, n_528;
  wire n_535, n_557, n_574, n_576, n_578, n_579, n_580, n_581;
  wire n_583, n_584, n_585, n_586, n_587, n_589, n_590, n_593;
  wire n_595, n_598, n_603, n_610, n_620, n_624, n_639, n_642;
  wire n_644, n_645, n_646, n_647, n_649, n_650, n_651, n_652;
  wire n_653, n_655, n_656, n_659, n_661, n_664, n_671, n_678;
  wire n_690, n_694, n_713, n_715, n_716, n_717, n_718, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_727, n_730, n_732;
  wire n_735, n_743, n_750, n_765, n_769, n_789, n_791, n_793;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_802;
  wire n_804, n_805, n_806, n_807, n_808, n_810, n_811, n_814;
  wire n_816, n_817, n_818, n_820, n_822, n_827, n_830, n_835;
  wire n_839, n_846, n_850, n_852, n_855, n_868, n_871, n_873;
  wire n_874, n_875, n_876, n_878, n_879, n_880, n_881, n_882;
  wire n_884, n_885, n_886, n_887, n_888, n_890, n_891, n_894;
  wire n_896, n_897, n_898, n_900, n_902, n_909, n_912, n_917;
  wire n_921, n_930, n_934, n_936, n_939, n_956, n_958, n_959;
  wire n_960, n_961, n_963, n_964, n_965, n_966, n_967, n_969;
  wire n_970, n_971, n_972, n_973, n_975, n_976, n_979, n_981;
  wire n_982, n_983, n_985, n_987, n_995, n_998, n_1003, n_1007;
  wire n_1019, n_1023, n_1025, n_1028, n_1045, n_1047, n_1052, n_1054;
  wire n_1058, n_1060, n_1064, n_1066, n_1070, n_1072, n_1075, n_1078;
  wire n_1080, n_1084, n_1086, n_1091, n_1099, n_1103, n_1106, n_1108;
  wire n_1146, n_1148, n_1152, n_1154, n_1158, n_1160, n_1164, n_1166;
  wire n_1169, n_1172, n_1174, n_1178, n_1180, n_1186, n_1187, n_1189;
  wire n_1197, n_1201, n_1247, n_1249, n_1253, n_1255, n_1259, n_1261;
  wire n_1265, n_1267, n_1270, n_1273, n_1275, n_1279, n_1281, n_1288;
  wire n_1293, n_1301, n_1305, n_1312, n_1342, n_1343, n_1344, n_1345;
  wire n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353;
  wire n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361;
  wire n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369;
  wire n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377;
  wire n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385;
  wire n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393;
  wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
  wire n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409;
  wire n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418;
  wire n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1427;
  wire n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435;
  wire n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443;
  wire n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468;
  wire n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484;
  wire n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508;
  wire n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517;
  wire n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525;
  wire n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557;
  wire n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565;
  wire n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572;
  nand g8 (QUOTIENT[9], n_46, n_49);
  nand g20 (QUOTIENT[7], n_66, n_69);
  nand g32 (QUOTIENT[5], n_94, n_97);
  nand g44 (QUOTIENT[3], n_132, n_135);
  or g55 (QUOTIENT[0], n_186, n_1572);
  xor g57 (n_277, B[0], B[1]);
  nand g58 (n_198, B[0], B[1]);
  nand g63 (n_204, B[1], B[2]);
  nand g9 (n_206, B[2], B[3]);
  nand g11 (n_208, B[3], B[4]);
  nand g65 (n_212, B[4], B[5]);
  nand g67 (n_214, B[5], B[6]);
  nand g69 (n_218, B[6], B[7]);
  nand g71 (n_220, B[7], B[8]);
  nand g21 (n_224, B[8], B[9]);
  nand g74 (n_228, n_204, n_1358);
  nor g75 (n_209, n_206, n_207);
  nor g78 (n_231, n_289, n_207);
  nor g79 (n_215, n_212, n_213);
  nor g34 (n_237, n_291, n_213);
  nor g35 (n_221, n_218, n_219);
  nor g82 (n_239, n_223, n_219);
  nand g45 (n_264, n_206, n_1390);
  nand g46 (n_233, n_231, n_228);
  nand g47 (n_244, n_1362, n_233);
  nor g48 (n_235, n_223, n_234);
  nand g95 (n_252, n_237, n_239);
  nand g98 (n_268, n_212, n_1402);
  nand g99 (n_247, n_237, n_244);
  nand g100 (n_270, n_234, n_247);
  nand g103 (n_273, n_1391, n_1403);
  nand g106 (n_256, n_1392, n_1404);
  nand g109 (n_276, n_224, n_1406);
  nand g110 (n_260, n_1345, n_256);
  xnor g115 (n_32, n_228, n_1359);
  xnor g118 (n_33, n_264, n_1361);
  xnor g120 (n_34, n_244, n_1363);
  xnor g123 (n_35, n_268, n_1364);
  xnor g125 (n_36, n_270, n_1365);
  xnor g128 (n_37, n_273, n_1367);
  xnor g130 (n_38, n_256, n_1369);
  nand g143 (n_286, n_284, n_1375);
  nor g144 (n_289, B[2], B[3]);
  nor g145 (n_291, B[4], B[5]);
  nor g146 (n_223, B[6], B[7]);
  nor g147 (n_307, B[8], B[9]);
  nand g150 (n_290, n_289, n_286);
  nand g153 (n_301, n_291, n_223);
  xnor g165 (n_42, n_282, n_1377);
  nand g191 (n_323, n_321, n_318);
  nor g192 (n_326, B[1], B[2]);
  nor g193 (n_207, B[3], B[4]);
  nor g194 (n_213, B[5], B[6]);
  nor g195 (n_219, B[7], B[8]);
  nand g198 (n_327, n_326, n_323);
  nand g201 (n_340, n_207, n_213);
  nand g245 (n_365, n_363, n_1389);
  nor g246 (n_368, n_31, n_32);
  nor g247 (n_370, n_33, n_34);
  nor g248 (n_372, n_35, n_36);
  nor g249 (n_373, n_37, n_38);
  nor g250 (n_375, n_1408, n_1407);
  nand g253 (n_369, n_368, n_365);
  nand g256 (n_383, n_370, n_372);
  nand g259 (n_393, n_373, n_375);
  xnor g275 (n_43, n_282, n_1393);
  nand g312 (n_420, n_412, n_1379);
  nor g313 (n_417, n_414, n_415);
  nor g316 (n_423, n_419, n_415);
  nand g322 (n_446, n_414, n_1417);
  nand g323 (n_425, n_423, n_420);
  nand g324 (n_429, n_1411, n_425);
  xnor g339 (n_56, n_410, n_1380);
  xnor g341 (n_58, n_420, n_1414);
  xnor g344 (n_61, n_446, n_1418);
  nand g371 (n_469, n_461, n_458);
  nor g372 (n_466, n_463, n_464);
  nor g375 (n_472, n_468, n_464);
  nand g381 (n_499, n_463, n_1419);
  nand g382 (n_474, n_472, n_469);
  nand g383 (n_480, n_1412, n_474);
  xnor g404 (n_59, n_469, n_1415);
  xnor g407 (n_62, n_499, n_1420);
  nand g437 (n_523, n_515, n_1394);
  nor g438 (n_520, n_517, n_518);
  nor g441 (n_526, n_522, n_518);
  nand g448 (n_557, n_517, n_1421);
  nand g449 (n_528, n_526, n_523);
  nand g450 (n_535, n_1413, n_528);
  xnor g472 (n_57, n_410, n_1395);
  xnor g474 (n_60, n_523, n_1416);
  xnor g477 (n_63, n_557, n_1422);
  nand g519 (n_590, n_576, n_1382);
  nor g520 (n_581, n_578, n_579);
  nor g523 (n_593, n_583, n_579);
  nor g524 (n_587, n_584, n_585);
  nor g527 (n_598, n_589, n_585);
  nand g532 (n_620, n_578, n_1436);
  nand g533 (n_595, n_593, n_590);
  nand g534 (n_603, n_1428, n_595);
  nand g540 (n_610, n_598, n_223);
  nand g543 (n_624, n_584, n_1454);
  nand g554 (n_92, n_307, n_1457);
  xnor g556 (n_78, n_574, n_1383);
  xnor g558 (n_80, n_590, n_1433);
  xnor g561 (n_83, n_620, n_1437);
  xnor g563 (n_86, n_603, n_1442);
  xnor g566 (n_89, n_624, n_1445);
  nand g596 (n_656, n_642, n_639);
  nor g597 (n_647, n_644, n_645);
  nor g600 (n_659, n_649, n_645);
  nor g601 (n_653, n_650, n_651);
  nor g604 (n_664, n_655, n_651);
  nand g609 (n_690, n_644, n_1438);
  nand g610 (n_661, n_659, n_656);
  nand g611 (n_671, n_1430, n_661);
  nand g617 (n_678, n_664, n_213);
  nand g622 (n_694, n_650, n_1455);
  xnor g639 (n_81, n_656, n_1434);
  xnor g642 (n_84, n_690, n_1439);
  xnor g644 (n_87, n_671, n_1443);
  xnor g647 (n_90, n_694, n_1446);
  nand g679 (n_727, n_713, n_1396);
  nor g680 (n_718, n_715, n_716);
  nor g683 (n_730, n_720, n_716);
  nor g684 (n_724, n_721, n_722);
  nor g687 (n_735, n_726, n_722);
  nand g693 (n_765, n_715, n_1440);
  nand g694 (n_732, n_730, n_727);
  nand g695 (n_743, n_1432, n_732);
  nand g701 (n_750, n_735, n_372);
  nand g707 (n_769, n_721, n_1456);
  xnor g724 (n_79, n_574, n_1397);
  xnor g726 (n_82, n_727, n_1435);
  xnor g729 (n_85, n_765, n_1441);
  xnor g731 (n_88, n_743, n_1444);
  xnor g734 (n_91, n_769, n_1447);
  nand g780 (n_811, n_791, n_1385);
  nor g781 (n_796, n_793, n_794);
  nor g784 (n_814, n_798, n_794);
  nor g785 (n_802, n_799, n_800);
  nor g788 (n_820, n_804, n_800);
  nor g789 (n_808, n_805, n_806);
  nor g792 (n_822, n_810, n_806);
  nand g796 (n_846, n_793, n_1479);
  nand g797 (n_816, n_814, n_811);
  nand g798 (n_827, n_1462, n_816);
  nor g799 (n_818, n_810, n_817);
  nand g808 (n_835, n_820, n_822);
  nand g811 (n_850, n_799, n_1506);
  nand g812 (n_830, n_820, n_827);
  nand g813 (n_852, n_817, n_830);
  nand g816 (n_855, n_1500, n_1501);
  nand g819 (n_839, n_1494, n_1495);
  nand g822 (n_130, n_307, n_839);
  xnor g824 (n_109, n_789, n_1386);
  xnor g826 (n_112, n_811, n_1476);
  xnor g829 (n_115, n_846, n_1480);
  xnor g831 (n_118, n_827, n_1485);
  xnor g834 (n_121, n_850, n_1488);
  xnor g836 (n_124, n_852, n_1467);
  xnor g839 (n_127, n_855, n_1471);
  nand g871 (n_891, n_871, n_868);
  nor g872 (n_876, n_873, n_874);
  nor g875 (n_894, n_878, n_874);
  nor g876 (n_882, n_879, n_880);
  nor g879 (n_900, n_884, n_880);
  nor g880 (n_888, n_885, n_886);
  nor g883 (n_902, n_890, n_886);
  nand g887 (n_930, n_873, n_1481);
  nand g888 (n_896, n_894, n_891);
  nand g889 (n_909, n_1464, n_896);
  nor g890 (n_898, n_890, n_897);
  nand g899 (n_917, n_900, n_902);
  nand g904 (n_934, n_879, n_1507);
  nand g905 (n_912, n_900, n_909);
  nand g906 (n_936, n_897, n_912);
  nand g909 (n_939, n_1502, n_1503);
  nand g912 (n_921, n_1496, n_1497);
  xnor g921 (n_113, n_891, n_1477);
  xnor g924 (n_116, n_930, n_1482);
  xnor g926 (n_119, n_909, n_1486);
  xnor g929 (n_122, n_934, n_1489);
  xnor g931 (n_125, n_936, n_1468);
  xnor g934 (n_128, n_939, n_1473);
  nand g968 (n_976, n_956, n_1398);
  nor g969 (n_961, n_958, n_959);
  nor g972 (n_979, n_963, n_959);
  nor g973 (n_967, n_964, n_965);
  nor g976 (n_985, n_969, n_965);
  nor g977 (n_973, n_970, n_971);
  nor g980 (n_987, n_975, n_971);
  nand g985 (n_1019, n_958, n_1483);
  nand g986 (n_981, n_979, n_976);
  nand g987 (n_995, n_1466, n_981);
  nor g988 (n_983, n_975, n_982);
  nand g997 (n_1003, n_985, n_987);
  nand g1003 (n_1023, n_964, n_1508);
  nand g1004 (n_998, n_985, n_995);
  nand g1005 (n_1025, n_982, n_998);
  nand g1008 (n_1028, n_1504, n_1505);
  nand g1011 (n_1007, n_1498, n_1499);
  xnor g1020 (n_111, n_789, n_1399);
  xnor g1022 (n_114, n_976, n_1478);
  xnor g1025 (n_117, n_1019, n_1484);
  xnor g1027 (n_120, n_995, n_1487);
  xnor g1030 (n_123, n_1023, n_1490);
  xnor g1032 (n_126, n_1025, n_1469);
  xnor g1035 (n_129, n_1028, n_1475);
  nand g1086 (n_1075, n_1355, n_1388);
  nor g1087 (n_1054, n_1530, n_1052);
  nor g1090 (n_1078, n_1532, n_1052);
  nor g1091 (n_1060, n_1525, n_1058);
  nor g1094 (n_1084, n_1533, n_1058);
  nor g1095 (n_1066, n_1528, n_1064);
  nor g1098 (n_1086, n_1527, n_1064);
  nor g1099 (n_1072, n_1522, n_1070);
  nor g1102 (n_1106, n_1524, n_1070);
  nand g1106 (n_1080, n_1078, n_1075);
  nand g1107 (n_1091, n_1554, n_1080);
  nand g1117 (n_1099, n_1084, n_1086);
  nand g1128 (n_1103, n_1565, n_1566);
  nand g1132 (n_1108, n_1106, n_1103);
  nand g1133 (n_1045, n_1551, n_1108);
  nand g1191 (n_1169, n_1353, n_1354);
  nor g1192 (n_1148, n_1517, n_1146);
  nor g1195 (n_1172, n_1519, n_1146);
  nor g1196 (n_1154, n_1512, n_1152);
  nor g1199 (n_1178, n_1520, n_1152);
  nor g1200 (n_1160, n_1515, n_1158);
  nor g1203 (n_1180, n_1514, n_1158);
  nor g1204 (n_1166, n_1510, n_1164);
  nor g1207 (n_1187, n_1521, n_1164);
  nand g1211 (n_1174, n_1172, n_1169);
  nand g1212 (n_1189, n_1549, n_1174);
  nand g1222 (n_1197, n_1178, n_1180);
  nor g1223 (n_1186, B[9], n_1546);
  nand g1236 (n_1201, n_1563, n_1564);
  nand g1304 (n_1270, n_1373, n_1400);
  nor g1305 (n_1249, n_1541, n_1247);
  nor g1308 (n_1273, n_1543, n_1247);
  nor g1309 (n_1255, n_1536, n_1253);
  nor g1312 (n_1279, n_1544, n_1253);
  nor g1313 (n_1261, n_1539, n_1259);
  nor g1316 (n_1281, n_1538, n_1259);
  nor g1317 (n_1267, n_1534, n_1265);
  nor g1320 (n_1288, n_1545, n_1265);
  nand g1325 (n_1275, n_1273, n_1270);
  nand g1326 (n_1293, n_1558, n_1275);
  nand g1336 (n_1301, n_1279, n_1281);
  nand g1342 (n_1312, n_1288, n_375);
  nand g1353 (n_1305, n_1567, n_1568);
  or g1404 (n_284, B[1], wc);
  not gc (wc, A[9]);
  or g1405 (n_282, wc0, A[8]);
  not gc0 (wc0, B[0]);
  and g1406 (n_1342, B[1], wc1);
  not gc1 (wc1, A[9]);
  or g1407 (n_321, B[0], wc2);
  not gc2 (wc2, A[9]);
  and g1408 (n_318, B[0], wc3);
  not gc3 (wc3, A[9]);
  or g1409 (n_1343, B[9], wc4);
  not gc4 (wc4, n_219);
  and g1410 (n_1344, B[9], wc5);
  not gc5 (wc5, n_224);
  and g1411 (n_1345, B[9], wc6);
  not gc6 (wc6, n_307);
  xnor g1412 (n_1346, A[8], B[0]);
  or g1413 (n_412, B[1], wc7);
  not gc7 (wc7, A[7]);
  or g1414 (n_410, wc8, A[6]);
  not gc8 (wc8, B[0]);
  and g1415 (n_1347, B[1], wc9);
  not gc9 (wc9, A[7]);
  or g1416 (n_461, B[0], wc10);
  not gc10 (wc10, A[7]);
  and g1417 (n_458, B[0], wc11);
  not gc11 (wc11, A[7]);
  xnor g1418 (n_1348, A[6], B[0]);
  or g1419 (n_576, B[1], wc12);
  not gc12 (wc12, A[5]);
  or g1420 (n_574, wc13, A[4]);
  not gc13 (wc13, B[0]);
  and g1421 (n_1349, B[1], wc14);
  not gc14 (wc14, A[5]);
  or g1422 (n_642, B[0], wc15);
  not gc15 (wc15, A[5]);
  and g1423 (n_639, B[0], wc16);
  not gc16 (wc16, A[5]);
  xnor g1424 (n_1350, A[4], B[0]);
  or g1425 (n_791, B[1], wc17);
  not gc17 (wc17, A[3]);
  or g1426 (n_789, wc18, A[2]);
  not gc18 (wc18, B[0]);
  and g1427 (n_1351, B[1], wc19);
  not gc19 (wc19, A[3]);
  or g1428 (n_871, B[0], wc20);
  not gc20 (wc20, A[3]);
  and g1429 (n_868, B[0], wc21);
  not gc21 (wc21, A[3]);
  xnor g1430 (n_1352, A[2], B[0]);
  or g1431 (n_1353, B[0], wc22);
  not gc22 (wc22, A[1]);
  and g1432 (n_1354, B[0], wc23);
  not gc23 (wc23, A[1]);
  or g1433 (n_1355, B[1], wc24);
  not gc24 (wc24, A[1]);
  or g1434 (n_1047, wc25, A[0]);
  not gc25 (wc25, B[0]);
  and g1435 (n_1356, B[1], wc26);
  not gc26 (wc26, A[1]);
  or g1436 (n_1357, n_326, wc27);
  not gc27 (wc27, n_204);
  or g1437 (n_1358, n_198, n_326);
  or g1438 (n_1359, n_289, wc28);
  not gc28 (wc28, n_206);
  or g1439 (n_363, wc29, n_277);
  not gc29 (wc29, A[9]);
  and g1440 (n_1360, wc30, n_277);
  not gc30 (wc30, A[9]);
  or g1441 (n_1361, n_207, wc31);
  not gc31 (wc31, n_208);
  and g1442 (n_1362, wc32, n_208);
  not gc32 (wc32, n_209);
  or g1443 (n_1363, n_291, wc33);
  not gc33 (wc33, n_212);
  or g1444 (n_1364, n_213, wc34);
  not gc34 (wc34, n_214);
  and g1445 (n_234, wc35, n_214);
  not gc35 (wc35, n_215);
  or g1446 (n_1365, n_223, wc36);
  not gc36 (wc36, n_218);
  or g1447 (n_1366, n_223, wc37);
  not gc37 (wc37, n_237);
  or g1448 (n_1367, n_219, wc38);
  not gc38 (wc38, n_220);
  and g1449 (n_1368, wc39, n_220);
  not gc39 (wc39, n_221);
  or g1450 (n_1369, n_307, wc40);
  not gc40 (wc40, n_224);
  or g1451 (n_515, wc41, n_277);
  not gc41 (wc41, A[7]);
  and g1452 (n_1370, wc42, n_277);
  not gc42 (wc42, A[7]);
  or g1453 (n_713, wc43, n_277);
  not gc43 (wc43, A[5]);
  and g1454 (n_1371, wc44, n_277);
  not gc44 (wc44, A[5]);
  or g1455 (n_956, wc45, n_277);
  not gc45 (wc45, A[3]);
  and g1456 (n_1372, wc46, n_277);
  not gc46 (wc46, A[3]);
  or g1457 (n_1373, wc47, n_277);
  not gc47 (wc47, A[1]);
  and g1458 (n_1374, wc48, n_277);
  not gc48 (wc48, A[1]);
  or g1459 (n_1375, n_1342, wc49);
  not gc49 (wc49, n_282);
  xor g1460 (n_31, n_198, n_1357);
  and g1461 (n_1376, wc50, n_239);
  not gc50 (wc50, n_234);
  or g1462 (n_1377, n_1342, wc51);
  not gc51 (wc51, n_284);
  or g1463 (n_1378, n_318, wc52);
  not gc52 (wc52, n_321);
  or g1464 (n_1379, n_1347, wc53);
  not gc53 (wc53, n_410);
  or g1465 (n_1380, n_1347, wc54);
  not gc54 (wc54, n_412);
  or g1466 (n_1381, n_458, wc55);
  not gc55 (wc55, n_461);
  or g1467 (n_1382, n_1349, wc56);
  not gc56 (wc56, n_574);
  or g1468 (n_1383, n_1349, wc57);
  not gc57 (wc57, n_576);
  or g1469 (n_1384, n_639, wc58);
  not gc58 (wc58, n_642);
  or g1470 (n_1385, n_1351, wc59);
  not gc59 (wc59, n_789);
  or g1471 (n_1386, n_1351, wc60);
  not gc60 (wc60, n_791);
  or g1472 (n_1387, n_868, wc61);
  not gc61 (wc61, n_871);
  or g1473 (n_1388, n_1356, wc62);
  not gc62 (wc62, n_1047);
  or g1474 (n_1389, n_1360, wc63);
  not gc63 (wc63, n_282);
  or g1475 (n_1390, n_289, wc64);
  not gc64 (wc64, n_228);
  and g1476 (n_1391, wc65, n_218);
  not gc65 (wc65, n_235);
  and g1477 (n_1392, wc66, n_1368);
  not gc66 (wc66, n_1376);
  or g1478 (n_1393, n_1360, wc67);
  not gc67 (wc67, n_363);
  or g1479 (n_1394, n_1370, wc68);
  not gc68 (wc68, n_410);
  or g1480 (n_1395, n_1370, wc69);
  not gc69 (wc69, n_515);
  or g1481 (n_1396, n_1371, wc70);
  not gc70 (wc70, n_574);
  or g1482 (n_1397, n_1371, wc71);
  not gc71 (wc71, n_713);
  or g1483 (n_1398, n_1372, wc72);
  not gc72 (wc72, n_789);
  or g1484 (n_1399, n_1372, wc73);
  not gc73 (wc73, n_956);
  or g1485 (n_1400, n_1374, wc74);
  not gc74 (wc74, n_1047);
  or g1486 (n_1401, n_327, n_340);
  or g1487 (n_1402, n_291, wc75);
  not gc75 (wc75, n_244);
  or g1488 (n_1403, n_1366, wc76);
  not gc76 (wc76, n_244);
  or g1489 (n_1404, n_252, wc77);
  not gc77 (wc77, n_244);
  or g1490 (n_1405, n_290, n_301);
  or g1491 (n_46, n_1343, n_1401);
  or g1492 (n_1406, n_307, wc78);
  not gc78 (wc78, n_256);
  or g1493 (n_44, n_1405, wc79);
  not gc79 (wc79, n_307);
  or g1494 (n_1407, n_1344, wc80);
  not gc80 (wc80, n_260);
  xor g1495 (n_1408, n_276, B[9]);
  and g1496 (n_47, wc81, n_46);
  not gc81 (wc81, n_44);
  or g1497 (n_1409, n_369, n_383);
  or g1498 (n_49, n_393, n_1409);
  and g1499 (n_50, n_49, wc82);
  not gc82 (wc82, n_46);
  or g1500 (QUOTIENT[8], wc83, n_47);
  not gc83 (wc83, n_49);
  or g1501 (n_53, wc84, wc85, wc87, wc88);
  and gc90 (wc88, wc89, wc90);
  not gc89 (wc90, n_1346);
  not gc88 (wc89, n_49);
  and gc87 (wc87, A[8], n_50);
  and gc86 (wc85, n_47, wc86);
  not gc85 (wc86, n_1346);
  and gc84 (wc84, A[8], n_44);
  or g1502 (n_54, wc91, wc92, wc93, wc94);
  and gc95 (wc94, wc95, n_43);
  not gc94 (wc95, n_49);
  and gc93 (wc93, n_50, n_1378);
  and gc92 (wc92, n_47, n_42);
  and gc91 (wc91, A[9], n_44);
  or g1503 (n_414, B[2], wc96);
  not gc96 (wc96, n_53);
  and g1504 (n_415, B[3], wc97);
  not gc97 (wc97, n_54);
  or g1505 (n_416, B[3], wc98);
  not gc98 (wc98, n_54);
  and g1506 (n_419, B[2], wc99);
  not gc99 (wc99, n_53);
  or g1507 (n_463, B[1], wc100);
  not gc100 (wc100, n_53);
  and g1508 (n_464, B[2], wc101);
  not gc101 (wc101, n_54);
  or g1509 (n_465, B[2], wc102);
  not gc102 (wc102, n_54);
  and g1510 (n_468, B[1], wc103);
  not gc103 (wc103, n_53);
  or g1511 (n_517, wc104, n_31);
  not gc104 (wc104, n_53);
  and g1512 (n_518, wc105, n_32);
  not gc105 (wc105, n_54);
  or g1513 (n_519, wc106, n_32);
  not gc106 (wc106, n_54);
  and g1514 (n_522, wc107, n_31);
  not gc107 (wc107, n_53);
  and g1515 (n_1411, n_416, wc108);
  not gc108 (wc108, n_417);
  and g1516 (n_1412, n_465, wc109);
  not gc109 (wc109, n_466);
  and g1517 (n_1413, n_519, wc110);
  not gc110 (wc110, n_520);
  or g1518 (n_1414, n_419, wc111);
  not gc111 (wc111, n_414);
  or g1519 (n_1415, n_468, wc112);
  not gc112 (wc112, n_463);
  or g1520 (n_1416, n_522, wc113);
  not gc113 (wc113, n_517);
  or g1521 (n_1417, n_419, wc114);
  not gc114 (wc114, n_420);
  or g1522 (n_1418, wc115, n_415);
  not gc115 (wc115, n_416);
  or g1523 (n_1419, n_468, wc116);
  not gc116 (wc116, n_469);
  or g1524 (n_1420, wc117, n_464);
  not gc117 (wc117, n_465);
  or g1525 (n_1421, n_522, wc118);
  not gc118 (wc118, n_523);
  or g1526 (n_1422, wc119, n_518);
  not gc119 (wc119, n_519);
  or g1527 (n_1423, wc120, n_301);
  not gc120 (wc120, n_429);
  or g1528 (n_1424, wc121, n_340);
  not gc121 (wc121, n_480);
  or g1529 (n_1425, wc122, n_383);
  not gc122 (wc122, n_535);
  or g1530 (n_64, n_1423, wc123);
  not gc123 (wc123, n_307);
  or g1531 (n_66, n_1343, n_1424);
  or g1532 (n_69, n_393, n_1425);
  and g1533 (n_67, n_66, wc124);
  not gc124 (wc124, n_64);
  and g1534 (n_70, n_69, wc125);
  not gc125 (wc125, n_66);
  or g1535 (QUOTIENT[6], n_67, wc126);
  not gc126 (wc126, n_69);
  or g1536 (n_75, wc127, wc128, wc129, wc130);
  and gc131 (wc130, wc131, n_60);
  not gc130 (wc131, n_69);
  and gc129 (wc129, n_70, n_59);
  and gc128 (wc128, n_67, n_58);
  and gc127 (wc127, n_64, n_53);
  or g1537 (n_76, wc132, wc133, wc134, wc135);
  and gc136 (wc135, wc136, n_63);
  not gc135 (wc136, n_69);
  and gc134 (wc134, n_70, n_62);
  and gc133 (wc133, n_67, n_61);
  and gc132 (wc132, n_64, n_54);
  or g1538 (n_73, wc137, wc138, wc140, wc141);
  and gc143 (wc141, wc142, wc143);
  not gc142 (wc143, n_1348);
  not gc141 (wc142, n_69);
  and gc140 (wc140, A[6], n_70);
  and gc139 (wc138, n_67, wc139);
  not gc138 (wc139, n_1348);
  and gc137 (wc137, A[6], n_64);
  or g1539 (n_74, wc144, wc145, wc146, wc147);
  and gc148 (wc147, wc148, n_57);
  not gc147 (wc148, n_69);
  and gc146 (wc146, n_70, n_1381);
  and gc145 (wc145, n_67, n_56);
  and gc144 (wc144, A[7], n_64);
  or g1540 (n_584, B[4], wc149);
  not gc149 (wc149, n_75);
  and g1541 (n_585, B[5], wc150);
  not gc150 (wc150, n_76);
  or g1542 (n_586, B[5], wc151);
  not gc151 (wc151, n_76);
  or g1543 (n_578, B[2], wc152);
  not gc152 (wc152, n_73);
  and g1544 (n_579, B[3], wc153);
  not gc153 (wc153, n_74);
  or g1545 (n_580, B[3], wc154);
  not gc154 (wc154, n_74);
  and g1546 (n_583, B[2], wc155);
  not gc155 (wc155, n_73);
  and g1547 (n_589, B[4], wc156);
  not gc156 (wc156, n_75);
  or g1548 (n_650, B[3], wc157);
  not gc157 (wc157, n_75);
  and g1549 (n_651, B[4], wc158);
  not gc158 (wc158, n_76);
  or g1550 (n_652, B[4], wc159);
  not gc159 (wc159, n_76);
  or g1551 (n_644, B[1], wc160);
  not gc160 (wc160, n_73);
  and g1552 (n_645, B[2], wc161);
  not gc161 (wc161, n_74);
  or g1553 (n_646, B[2], wc162);
  not gc162 (wc162, n_74);
  and g1554 (n_649, B[1], wc163);
  not gc163 (wc163, n_73);
  and g1555 (n_655, B[3], wc164);
  not gc164 (wc164, n_75);
  or g1556 (n_721, wc165, n_33);
  not gc165 (wc165, n_75);
  and g1557 (n_722, wc166, n_34);
  not gc166 (wc166, n_76);
  or g1558 (n_723, wc167, n_34);
  not gc167 (wc167, n_76);
  or g1559 (n_715, wc168, n_31);
  not gc168 (wc168, n_73);
  and g1560 (n_716, wc169, n_32);
  not gc169 (wc169, n_74);
  or g1561 (n_717, wc170, n_32);
  not gc170 (wc170, n_74);
  and g1562 (n_720, wc171, n_31);
  not gc171 (wc171, n_73);
  and g1563 (n_726, wc172, n_33);
  not gc172 (wc172, n_75);
  and g1564 (n_1427, n_586, wc173);
  not gc173 (wc173, n_587);
  and g1565 (n_1428, n_580, wc174);
  not gc174 (wc174, n_581);
  and g1566 (n_1429, n_652, wc175);
  not gc175 (wc175, n_653);
  and g1567 (n_1430, n_646, wc176);
  not gc176 (wc176, n_647);
  and g1568 (n_1431, n_723, wc177);
  not gc177 (wc177, n_724);
  and g1569 (n_1432, n_717, wc178);
  not gc178 (wc178, n_718);
  or g1570 (n_1433, n_583, wc179);
  not gc179 (wc179, n_578);
  or g1571 (n_1434, n_649, wc180);
  not gc180 (wc180, n_644);
  or g1572 (n_1435, n_720, wc181);
  not gc181 (wc181, n_715);
  or g1573 (n_1436, n_583, wc182);
  not gc182 (wc182, n_590);
  or g1574 (n_1437, wc183, n_579);
  not gc183 (wc183, n_580);
  or g1575 (n_1438, n_649, wc184);
  not gc184 (wc184, n_656);
  or g1576 (n_1439, wc185, n_645);
  not gc185 (wc185, n_646);
  or g1577 (n_1440, n_720, wc186);
  not gc186 (wc186, n_727);
  or g1578 (n_1441, wc187, n_716);
  not gc187 (wc187, n_717);
  or g1579 (n_1442, n_589, wc188);
  not gc188 (wc188, n_584);
  or g1580 (n_1443, n_655, wc189);
  not gc189 (wc189, n_650);
  or g1581 (n_1444, n_726, wc190);
  not gc190 (wc190, n_721);
  or g1582 (n_1445, wc191, n_585);
  not gc191 (wc191, n_586);
  or g1583 (n_1446, wc192, n_651);
  not gc192 (wc192, n_652);
  or g1584 (n_1447, wc193, n_722);
  not gc193 (wc193, n_723);
  and g1585 (n_1448, wc194, n_223);
  not gc194 (wc194, n_1427);
  and g1586 (n_1449, wc195, n_213);
  not gc195 (wc195, n_1429);
  and g1587 (n_1450, wc196, n_372);
  not gc196 (wc196, n_1431);
  or g1588 (n_1451, n_610, wc197);
  not gc197 (wc197, n_603);
  or g1589 (n_1452, n_678, wc198);
  not gc198 (wc198, n_671);
  or g1590 (n_1453, n_750, wc199);
  not gc199 (wc199, n_743);
  or g1591 (n_1454, n_589, wc200);
  not gc200 (wc200, n_603);
  or g1592 (n_1455, n_655, wc201);
  not gc201 (wc201, n_671);
  or g1593 (n_1456, n_726, wc202);
  not gc202 (wc202, n_743);
  or g1594 (n_1457, wc203, n_1448);
  not gc203 (wc203, n_1451);
  or g1595 (n_1458, wc204, n_1449);
  not gc204 (wc204, n_1452);
  or g1596 (n_1459, wc205, n_1450);
  not gc205 (wc205, n_1453);
  or g1597 (n_94, wc206, n_1343);
  not gc206 (wc206, n_1458);
  or g1598 (n_97, wc207, n_393);
  not gc207 (wc207, n_1459);
  and g1599 (n_95, n_94, wc208);
  not gc208 (wc208, n_92);
  and g1600 (n_98, n_97, wc209);
  not gc209 (wc209, n_94);
  or g1601 (QUOTIENT[4], n_95, wc210);
  not gc210 (wc210, n_97);
  or g1602 (n_103, wc211, wc212, wc213, wc214);
  and gc215 (wc214, wc215, n_82);
  not gc214 (wc215, n_97);
  and gc213 (wc213, n_98, n_81);
  and gc212 (wc212, n_95, n_80);
  and gc211 (wc211, n_73, n_92);
  or g1603 (n_104, wc216, wc217, wc218, wc219);
  and gc220 (wc219, wc220, n_85);
  not gc219 (wc220, n_97);
  and gc218 (wc218, n_98, n_84);
  and gc217 (wc217, n_95, n_83);
  and gc216 (wc216, n_74, n_92);
  or g1604 (n_105, wc221, wc222, wc223, wc224);
  and gc225 (wc224, wc225, n_88);
  not gc224 (wc225, n_97);
  and gc223 (wc223, n_98, n_87);
  and gc222 (wc222, n_95, n_86);
  and gc221 (wc221, n_75, n_92);
  or g1605 (n_106, wc226, wc227, wc228, wc229);
  and gc230 (wc229, wc230, n_91);
  not gc229 (wc230, n_97);
  and gc228 (wc228, n_98, n_90);
  and gc227 (wc227, n_95, n_89);
  and gc226 (wc226, n_76, n_92);
  or g1606 (n_101, wc231, wc232, wc234, wc235);
  and gc237 (wc235, wc236, wc237);
  not gc236 (wc237, n_1350);
  not gc235 (wc236, n_97);
  and gc234 (wc234, A[4], n_98);
  and gc233 (wc232, n_95, wc233);
  not gc232 (wc233, n_1350);
  and gc231 (wc231, A[4], n_92);
  or g1607 (n_102, wc238, wc239, wc240, wc241);
  and gc242 (wc241, wc242, n_79);
  not gc241 (wc242, n_97);
  and gc240 (wc240, n_98, n_1384);
  and gc239 (wc239, n_95, n_78);
  and gc238 (wc238, A[5], n_92);
  or g1608 (n_799, B[4], wc243);
  not gc243 (wc243, n_103);
  and g1609 (n_800, B[5], wc244);
  not gc244 (wc244, n_104);
  or g1610 (n_801, B[5], wc245);
  not gc245 (wc245, n_104);
  and g1611 (n_810, B[6], wc246);
  not gc246 (wc246, n_105);
  and g1612 (n_806, B[7], wc247);
  not gc247 (wc247, n_106);
  or g1613 (n_805, B[6], wc248);
  not gc248 (wc248, n_105);
  or g1614 (n_807, B[7], wc249);
  not gc249 (wc249, n_106);
  or g1615 (n_793, B[2], wc250);
  not gc250 (wc250, n_101);
  and g1616 (n_794, B[3], wc251);
  not gc251 (wc251, n_102);
  or g1617 (n_795, B[3], wc252);
  not gc252 (wc252, n_102);
  and g1618 (n_798, B[2], wc253);
  not gc253 (wc253, n_101);
  and g1619 (n_804, B[4], wc254);
  not gc254 (wc254, n_103);
  or g1620 (n_879, B[3], wc255);
  not gc255 (wc255, n_103);
  and g1621 (n_880, B[4], wc256);
  not gc256 (wc256, n_104);
  or g1622 (n_881, B[4], wc257);
  not gc257 (wc257, n_104);
  and g1623 (n_890, B[5], wc258);
  not gc258 (wc258, n_105);
  and g1624 (n_886, B[6], wc259);
  not gc259 (wc259, n_106);
  or g1625 (n_885, B[5], wc260);
  not gc260 (wc260, n_105);
  or g1626 (n_887, B[6], wc261);
  not gc261 (wc261, n_106);
  or g1627 (n_873, B[1], wc262);
  not gc262 (wc262, n_101);
  and g1628 (n_874, B[2], wc263);
  not gc263 (wc263, n_102);
  or g1629 (n_875, B[2], wc264);
  not gc264 (wc264, n_102);
  and g1630 (n_878, B[1], wc265);
  not gc265 (wc265, n_101);
  and g1631 (n_884, B[3], wc266);
  not gc266 (wc266, n_103);
  or g1632 (n_964, wc267, n_33);
  not gc267 (wc267, n_103);
  and g1633 (n_965, wc268, n_34);
  not gc268 (wc268, n_104);
  or g1634 (n_966, wc269, n_34);
  not gc269 (wc269, n_104);
  and g1635 (n_975, wc270, n_35);
  not gc270 (wc270, n_105);
  and g1636 (n_971, wc271, n_36);
  not gc271 (wc271, n_106);
  or g1637 (n_970, wc272, n_35);
  not gc272 (wc272, n_105);
  or g1638 (n_972, wc273, n_36);
  not gc273 (wc273, n_106);
  or g1639 (n_958, wc274, n_31);
  not gc274 (wc274, n_101);
  and g1640 (n_959, wc275, n_32);
  not gc275 (wc275, n_102);
  or g1641 (n_960, wc276, n_32);
  not gc276 (wc276, n_102);
  and g1642 (n_963, wc277, n_31);
  not gc277 (wc277, n_101);
  and g1643 (n_969, wc278, n_33);
  not gc278 (wc278, n_103);
  and g1644 (n_817, n_801, wc279);
  not gc279 (wc279, n_802);
  and g1645 (n_1461, n_807, wc280);
  not gc280 (wc280, n_808);
  and g1646 (n_1462, n_795, wc281);
  not gc281 (wc281, n_796);
  and g1647 (n_897, n_881, wc282);
  not gc282 (wc282, n_882);
  and g1648 (n_1463, n_887, wc283);
  not gc283 (wc283, n_888);
  and g1649 (n_1464, n_875, wc284);
  not gc284 (wc284, n_876);
  and g1650 (n_982, n_966, wc285);
  not gc285 (wc285, n_967);
  and g1651 (n_1465, n_972, wc286);
  not gc286 (wc286, n_973);
  and g1652 (n_1466, n_960, wc287);
  not gc287 (wc287, n_961);
  or g1653 (n_1467, wc288, n_810);
  not gc288 (wc288, n_805);
  or g1654 (n_1468, wc289, n_890);
  not gc289 (wc289, n_885);
  or g1655 (n_1469, wc290, n_975);
  not gc290 (wc290, n_970);
  or g1656 (n_1470, n_810, wc291);
  not gc291 (wc291, n_820);
  or g1657 (n_1471, wc292, n_806);
  not gc292 (wc292, n_807);
  or g1658 (n_1472, n_890, wc293);
  not gc293 (wc293, n_900);
  or g1659 (n_1473, wc294, n_886);
  not gc294 (wc294, n_887);
  or g1660 (n_1474, n_975, wc295);
  not gc295 (wc295, n_985);
  or g1661 (n_1475, wc296, n_971);
  not gc296 (wc296, n_972);
  or g1662 (n_1476, n_798, wc297);
  not gc297 (wc297, n_793);
  or g1663 (n_1477, n_878, wc298);
  not gc298 (wc298, n_873);
  or g1664 (n_1478, n_963, wc299);
  not gc299 (wc299, n_958);
  or g1665 (n_1479, n_798, wc300);
  not gc300 (wc300, n_811);
  or g1666 (n_1480, wc301, n_794);
  not gc301 (wc301, n_795);
  or g1667 (n_1481, n_878, wc302);
  not gc302 (wc302, n_891);
  or g1668 (n_1482, wc303, n_874);
  not gc303 (wc303, n_875);
  or g1669 (n_1483, n_963, wc304);
  not gc304 (wc304, n_976);
  or g1670 (n_1484, wc305, n_959);
  not gc305 (wc305, n_960);
  or g1671 (n_1485, n_804, wc306);
  not gc306 (wc306, n_799);
  or g1672 (n_1486, n_884, wc307);
  not gc307 (wc307, n_879);
  or g1673 (n_1487, n_969, wc308);
  not gc308 (wc308, n_964);
  or g1674 (n_1488, wc309, n_800);
  not gc309 (wc309, n_801);
  or g1675 (n_1489, wc310, n_880);
  not gc310 (wc310, n_881);
  or g1676 (n_1490, wc311, n_965);
  not gc311 (wc311, n_966);
  and g1677 (n_1491, wc312, n_822);
  not gc312 (wc312, n_817);
  and g1678 (n_1492, wc313, n_902);
  not gc313 (wc313, n_897);
  and g1679 (n_1493, wc314, n_987);
  not gc314 (wc314, n_982);
  and g1680 (n_1494, wc315, n_1461);
  not gc315 (wc315, n_1491);
  or g1681 (n_1495, n_835, wc316);
  not gc316 (wc316, n_827);
  and g1682 (n_1496, wc317, n_1463);
  not gc317 (wc317, n_1492);
  or g1683 (n_1497, n_917, wc318);
  not gc318 (wc318, n_909);
  and g1684 (n_1498, wc319, n_1465);
  not gc319 (wc319, n_1493);
  or g1685 (n_1499, n_1003, wc320);
  not gc320 (wc320, n_995);
  and g1686 (n_1500, n_805, wc321);
  not gc321 (wc321, n_818);
  or g1687 (n_1501, n_1470, wc322);
  not gc322 (wc322, n_827);
  and g1688 (n_1502, n_885, wc323);
  not gc323 (wc323, n_898);
  or g1689 (n_1503, n_1472, wc324);
  not gc324 (wc324, n_909);
  and g1690 (n_1504, n_970, wc325);
  not gc325 (wc325, n_983);
  or g1691 (n_1505, n_1474, wc326);
  not gc326 (wc326, n_995);
  or g1692 (n_1506, n_804, wc327);
  not gc327 (wc327, n_827);
  or g1693 (n_1507, n_884, wc328);
  not gc328 (wc328, n_909);
  or g1694 (n_1508, n_969, wc329);
  not gc329 (wc329, n_995);
  or g1695 (n_132, n_1343, wc330);
  not gc330 (wc330, n_921);
  or g1696 (n_135, wc331, n_393);
  not gc331 (wc331, n_1007);
  and g1697 (n_133, n_132, wc332);
  not gc332 (wc332, n_130);
  and g1698 (n_136, n_135, wc333);
  not gc333 (wc333, n_132);
  or g1699 (QUOTIENT[2], n_133, wc334);
  not gc334 (wc334, n_135);
  or g1700 (n_147, wc335, wc336, wc337, wc338);
  and gc339 (wc338, wc339, n_126);
  not gc338 (wc339, n_135);
  and gc337 (wc337, n_136, n_125);
  and gc336 (wc336, n_133, n_124);
  and gc335 (wc335, n_105, n_130);
  or g1701 (n_148, wc340, wc341, wc342, wc343);
  and gc344 (wc343, wc344, n_129);
  not gc343 (wc344, n_135);
  and gc342 (wc342, n_136, n_128);
  and gc341 (wc341, n_133, n_127);
  and gc340 (wc340, n_106, n_130);
  or g1702 (n_143, wc345, wc346, wc347, wc348);
  and gc349 (wc348, wc349, n_114);
  not gc348 (wc349, n_135);
  and gc347 (wc347, n_136, n_113);
  and gc346 (wc346, n_133, n_112);
  and gc345 (wc345, n_101, n_130);
  or g1703 (n_144, wc350, wc351, wc352, wc353);
  and gc354 (wc353, wc354, n_117);
  not gc353 (wc354, n_135);
  and gc352 (wc352, n_136, n_116);
  and gc351 (wc351, n_133, n_115);
  and gc350 (wc350, n_102, n_130);
  or g1704 (n_145, wc355, wc356, wc357, wc358);
  and gc359 (wc358, wc359, n_120);
  not gc358 (wc359, n_135);
  and gc357 (wc357, n_136, n_119);
  and gc356 (wc356, n_133, n_118);
  and gc355 (wc355, n_103, n_130);
  or g1705 (n_146, wc360, wc361, wc362, wc363);
  and gc364 (wc363, wc364, n_123);
  not gc363 (wc364, n_135);
  and gc362 (wc362, n_136, n_122);
  and gc361 (wc361, n_133, n_121);
  and gc360 (wc360, n_104, n_130);
  or g1706 (n_141, wc365, wc366, wc368, wc369);
  and gc371 (wc369, wc370, wc371);
  not gc370 (wc371, n_1352);
  not gc369 (wc370, n_135);
  and gc368 (wc368, A[2], n_136);
  and gc367 (wc366, n_133, wc367);
  not gc366 (wc367, n_1352);
  and gc365 (wc365, A[2], n_130);
  or g1707 (n_142, wc372, wc373, wc374, wc375);
  and gc376 (wc375, wc376, n_111);
  not gc375 (wc376, n_135);
  and gc374 (wc374, n_136, n_1387);
  and gc373 (wc373, n_133, n_109);
  and gc372 (wc372, A[3], n_130);
  or g1708 (n_1510, B[7], wc377);
  not gc377 (wc377, n_147);
  and g1709 (n_1164, B[8], wc378);
  not gc378 (wc378, n_148);
  or g1710 (n_1511, B[8], wc379);
  not gc379 (wc379, n_148);
  or g1711 (n_1512, B[3], wc380);
  not gc380 (wc380, n_143);
  and g1712 (n_1152, B[4], wc381);
  not gc381 (wc381, n_144);
  or g1713 (n_1513, B[4], wc382);
  not gc382 (wc382, n_144);
  and g1714 (n_1514, B[5], wc383);
  not gc383 (wc383, n_145);
  and g1715 (n_1158, B[6], wc384);
  not gc384 (wc384, n_146);
  or g1716 (n_1515, B[5], wc385);
  not gc385 (wc385, n_145);
  or g1717 (n_1516, B[6], wc386);
  not gc386 (wc386, n_146);
  or g1718 (n_1517, B[1], wc387);
  not gc387 (wc387, n_141);
  and g1719 (n_1146, B[2], wc388);
  not gc388 (wc388, n_142);
  or g1720 (n_1518, B[2], wc389);
  not gc389 (wc389, n_142);
  and g1721 (n_1519, B[1], wc390);
  not gc390 (wc390, n_141);
  and g1722 (n_1520, B[3], wc391);
  not gc391 (wc391, n_143);
  and g1723 (n_1521, B[7], wc392);
  not gc392 (wc392, n_147);
  or g1724 (n_1522, B[8], wc393);
  not gc393 (wc393, n_147);
  and g1725 (n_1070, B[9], wc394);
  not gc394 (wc394, n_148);
  or g1726 (n_1523, B[9], wc395);
  not gc395 (wc395, n_148);
  and g1727 (n_1524, B[8], wc396);
  not gc396 (wc396, n_147);
  or g1728 (n_1525, B[4], wc397);
  not gc397 (wc397, n_143);
  and g1729 (n_1058, B[5], wc398);
  not gc398 (wc398, n_144);
  or g1730 (n_1526, B[5], wc399);
  not gc399 (wc399, n_144);
  and g1731 (n_1527, B[6], wc400);
  not gc400 (wc400, n_145);
  and g1732 (n_1064, B[7], wc401);
  not gc401 (wc401, n_146);
  or g1733 (n_1528, B[6], wc402);
  not gc402 (wc402, n_145);
  or g1734 (n_1529, B[7], wc403);
  not gc403 (wc403, n_146);
  or g1735 (n_1530, B[2], wc404);
  not gc404 (wc404, n_141);
  and g1736 (n_1052, B[3], wc405);
  not gc405 (wc405, n_142);
  or g1737 (n_1531, B[3], wc406);
  not gc406 (wc406, n_142);
  and g1738 (n_1532, B[2], wc407);
  not gc407 (wc407, n_141);
  and g1739 (n_1533, B[4], wc408);
  not gc408 (wc408, n_143);
  or g1740 (n_1534, wc409, n_37);
  not gc409 (wc409, n_147);
  and g1741 (n_1265, wc410, n_38);
  not gc410 (wc410, n_148);
  or g1742 (n_1535, wc411, n_38);
  not gc411 (wc411, n_148);
  or g1743 (n_1536, wc412, n_33);
  not gc412 (wc412, n_143);
  and g1744 (n_1253, wc413, n_34);
  not gc413 (wc413, n_144);
  or g1745 (n_1537, wc414, n_34);
  not gc414 (wc414, n_144);
  and g1746 (n_1538, wc415, n_35);
  not gc415 (wc415, n_145);
  and g1747 (n_1259, wc416, n_36);
  not gc416 (wc416, n_146);
  or g1748 (n_1539, wc417, n_35);
  not gc417 (wc417, n_145);
  or g1749 (n_1540, wc418, n_36);
  not gc418 (wc418, n_146);
  or g1750 (n_1541, wc419, n_31);
  not gc419 (wc419, n_141);
  and g1751 (n_1247, wc420, n_32);
  not gc420 (wc420, n_142);
  or g1752 (n_1542, wc421, n_32);
  not gc421 (wc421, n_142);
  and g1753 (n_1543, wc422, n_31);
  not gc422 (wc422, n_141);
  and g1754 (n_1544, wc423, n_33);
  not gc423 (wc423, n_143);
  and g1755 (n_1545, wc424, n_37);
  not gc424 (wc424, n_147);
  and g1756 (n_1546, n_1511, wc425);
  not gc425 (wc425, n_1166);
  and g1757 (n_1547, n_1513, wc426);
  not gc426 (wc426, n_1154);
  and g1758 (n_1548, n_1516, wc427);
  not gc427 (wc427, n_1160);
  and g1759 (n_1549, n_1518, wc428);
  not gc428 (wc428, n_1148);
  or g1760 (n_1550, B[9], wc429);
  not gc429 (wc429, n_1187);
  and g1761 (n_1551, n_1523, wc430);
  not gc430 (wc430, n_1072);
  and g1762 (n_1552, n_1526, wc431);
  not gc431 (wc431, n_1060);
  and g1763 (n_1553, n_1529, wc432);
  not gc432 (wc432, n_1066);
  and g1764 (n_1554, n_1531, wc433);
  not gc433 (wc433, n_1054);
  and g1765 (n_1555, n_1535, wc434);
  not gc434 (wc434, n_1267);
  and g1766 (n_1556, n_1537, wc435);
  not gc435 (wc435, n_1255);
  and g1767 (n_1557, n_1540, wc436);
  not gc436 (wc436, n_1261);
  and g1768 (n_1558, n_1542, wc437);
  not gc437 (wc437, n_1249);
  and g1769 (n_1559, wc438, n_1180);
  not gc438 (wc438, n_1547);
  and g1770 (n_1560, wc439, n_1086);
  not gc439 (wc439, n_1552);
  and g1771 (n_1561, wc440, n_375);
  not gc440 (wc440, n_1555);
  and g1772 (n_1562, wc441, n_1281);
  not gc441 (wc441, n_1556);
  and g1773 (n_1563, wc442, n_1548);
  not gc442 (wc442, n_1559);
  or g1774 (n_1564, n_1197, wc443);
  not gc443 (wc443, n_1189);
  and g1775 (n_1565, wc444, n_1553);
  not gc444 (wc444, n_1560);
  or g1776 (n_1566, n_1099, wc445);
  not gc445 (wc445, n_1091);
  and g1777 (n_1567, wc446, n_1557);
  not gc446 (wc446, n_1562);
  or g1778 (n_1568, n_1301, wc447);
  not gc447 (wc447, n_1293);
  or g1779 (n_1569, n_1550, wc448);
  not gc448 (wc448, n_1201);
  or g1780 (n_1570, wc449, n_1312);
  not gc449 (wc449, n_1305);
  or g1781 (n_1571, wc450, n_1186);
  not gc450 (wc450, n_1569);
  or g1782 (n_186, wc451, n_1561);
  not gc451 (wc451, n_1570);
  and g1783 (n_1572, wc452, n_1045);
  not gc452 (wc452, n_1571);
  or g1784 (QUOTIENT[1], n_1571, n_186);
endmodule

module divide_unsigned_16_GENERIC(A, B, QUOTIENT);
  input [9:0] A, B;
  output [9:0] QUOTIENT;
  wire [9:0] A, B;
  wire [9:0] QUOTIENT;
  divide_unsigned_16_GENERIC_REAL g1(.A (A), .B (B), .QUOTIENT
       (QUOTIENT));
endmodule

