library verilog;
use verilog.vl_types.all;
entity TestFixture is
end TestFixture;
