library verilog;
use verilog.vl_types.all;
entity lab1_tb is
end lab1_tb;
