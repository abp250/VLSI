library verilog;
use verilog.vl_types.all;
entity ALT_MULTADD_pipe_tb is
end ALT_MULTADD_pipe_tb;
