module add_unsigned_108_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [16:0] A, B;
  output [16:0] Z;
  wire [16:0] A, B;
  wire [16:0] Z;
  wire n_53, n_58, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_136, n_142, n_143;
  nand g1 (n_53, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_58, A[1], B[1]);
  nand g10 (n_62, n_58, n_142, n_143);
  xor g11 (n_61, A[1], B[1]);
  nand g13 (n_63, A[2], B[2]);
  nand g14 (n_64, A[2], n_62);
  nand g15 (n_65, B[2], n_62);
  nand g16 (n_67, n_63, n_64, n_65);
  xor g17 (n_66, A[2], B[2]);
  xor g18 (Z[2], n_62, n_66);
  nand g19 (n_68, A[3], B[3]);
  nand g20 (n_69, A[3], n_67);
  nand g21 (n_70, B[3], n_67);
  nand g22 (n_72, n_68, n_69, n_70);
  xor g23 (n_71, A[3], B[3]);
  xor g24 (Z[3], n_67, n_71);
  nand g25 (n_73, A[4], B[4]);
  nand g26 (n_74, A[4], n_72);
  nand g27 (n_75, B[4], n_72);
  nand g28 (n_77, n_73, n_74, n_75);
  xor g29 (n_76, A[4], B[4]);
  xor g30 (Z[4], n_72, n_76);
  nand g31 (n_78, A[5], B[5]);
  nand g32 (n_79, A[5], n_77);
  nand g33 (n_80, B[5], n_77);
  nand g34 (n_82, n_78, n_79, n_80);
  xor g35 (n_81, A[5], B[5]);
  xor g36 (Z[5], n_77, n_81);
  nand g37 (n_83, A[6], B[6]);
  nand g38 (n_84, A[6], n_82);
  nand g39 (n_85, B[6], n_82);
  nand g40 (n_87, n_83, n_84, n_85);
  xor g41 (n_86, A[6], B[6]);
  xor g42 (Z[6], n_82, n_86);
  nand g43 (n_88, A[7], B[7]);
  nand g44 (n_89, A[7], n_87);
  nand g45 (n_90, B[7], n_87);
  nand g46 (n_92, n_88, n_89, n_90);
  xor g47 (n_91, A[7], B[7]);
  xor g48 (Z[7], n_87, n_91);
  nand g49 (n_93, A[8], B[8]);
  nand g50 (n_94, A[8], n_92);
  nand g51 (n_95, B[8], n_92);
  nand g52 (n_97, n_93, n_94, n_95);
  xor g53 (n_96, A[8], B[8]);
  xor g54 (Z[8], n_92, n_96);
  nand g55 (n_98, A[9], B[9]);
  nand g56 (n_99, A[9], n_97);
  nand g57 (n_100, B[9], n_97);
  nand g58 (n_102, n_98, n_99, n_100);
  xor g59 (n_101, A[9], B[9]);
  xor g60 (Z[9], n_97, n_101);
  nand g61 (n_103, A[10], B[10]);
  nand g62 (n_104, A[10], n_102);
  nand g63 (n_105, B[10], n_102);
  nand g64 (n_107, n_103, n_104, n_105);
  xor g65 (n_106, A[10], B[10]);
  xor g66 (Z[10], n_102, n_106);
  nand g67 (n_108, A[11], B[11]);
  nand g68 (n_109, A[11], n_107);
  nand g69 (n_110, B[11], n_107);
  nand g70 (n_112, n_108, n_109, n_110);
  xor g71 (n_111, A[11], B[11]);
  xor g72 (Z[11], n_107, n_111);
  nand g73 (n_113, A[12], B[12]);
  nand g74 (n_114, A[12], n_112);
  nand g75 (n_115, B[12], n_112);
  nand g76 (n_117, n_113, n_114, n_115);
  xor g77 (n_116, A[12], B[12]);
  xor g78 (Z[12], n_112, n_116);
  nand g79 (n_118, A[13], B[13]);
  nand g80 (n_119, A[13], n_117);
  nand g81 (n_120, B[13], n_117);
  nand g82 (n_122, n_118, n_119, n_120);
  xor g83 (n_121, A[13], B[13]);
  xor g84 (Z[13], n_117, n_121);
  nand g85 (n_123, A[14], B[14]);
  nand g86 (n_124, A[14], n_122);
  nand g87 (n_125, B[14], n_122);
  nand g88 (n_127, n_123, n_124, n_125);
  xor g89 (n_126, A[14], B[14]);
  xor g90 (Z[14], n_122, n_126);
  nand g91 (n_128, A[15], B[15]);
  nand g92 (n_129, A[15], n_127);
  nand g93 (n_130, B[15], n_127);
  nand g94 (n_132, n_128, n_129, n_130);
  xor g95 (n_131, A[15], B[15]);
  xor g96 (Z[15], n_127, n_131);
  xor g101 (n_136, A[16], B[16]);
  xor g102 (Z[16], n_132, n_136);
  or g104 (n_142, wc, n_53);
  not gc (wc, A[1]);
  or g105 (n_143, wc0, n_53);
  not gc0 (wc0, B[1]);
  xnor g106 (Z[1], n_53, n_61);
endmodule

module add_unsigned_108_GENERIC(A, B, Z);
  input [16:0] A, B;
  output [16:0] Z;
  wire [16:0] A, B;
  wire [16:0] Z;
  add_unsigned_108_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module csa_tree_GENERIC_REAL(in_0, in_1, in_2, in_3, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( in_0 * in_1 )  + ( in_2 * in_3 )  )  ; assign out_1 = 17'b0;"
  input [7:0] in_0, in_1, in_2, in_3;
  output [16:0] out_0, out_1;
  wire [7:0] in_0, in_1, in_2, in_3;
  wire [16:0] out_0, out_1;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697;
  wire n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  assign out_1[16] = 1'b0;
  assign out_0[16] = 1'b0;
  and g1 (out_0[0], in_0[0], in_1[0]);
  and g2 (n_33, in_0[1], in_1[0]);
  and g3 (n_36, in_0[2], in_1[0]);
  and g4 (n_44, in_0[3], in_1[0]);
  and g5 (n_58, in_0[4], in_1[0]);
  and g6 (n_78, in_0[5], in_1[0]);
  and g7 (n_104, in_0[6], in_1[0]);
  and g8 (n_136, in_0[7], in_1[0]);
  and g9 (out_0[1], in_0[0], in_1[1]);
  and g10 (n_37, in_0[1], in_1[1]);
  and g11 (n_45, in_0[2], in_1[1]);
  and g12 (n_59, in_0[3], in_1[1]);
  and g13 (n_79, in_0[4], in_1[1]);
  and g14 (n_105, in_0[5], in_1[1]);
  and g15 (n_137, in_0[6], in_1[1]);
  and g16 (n_174, in_0[7], in_1[1]);
  and g17 (n_41, in_0[0], in_1[2]);
  and g18 (n_49, in_0[1], in_1[2]);
  and g19 (n_65, in_0[2], in_1[2]);
  and g20 (n_86, in_0[3], in_1[2]);
  and g21 (n_112, in_0[4], in_1[2]);
  and g22 (n_145, in_0[5], in_1[2]);
  and g23 (n_175, in_0[6], in_1[2]);
  and g24 (n_212, in_0[7], in_1[2]);
  and g25 (n_46, in_0[0], in_1[3]);
  and g26 (n_60, in_0[1], in_1[3]);
  and g27 (n_80, in_0[2], in_1[3]);
  and g28 (n_106, in_0[3], in_1[3]);
  and g29 (n_138, in_0[4], in_1[3]);
  and g30 (n_182, in_0[5], in_1[3]);
  and g31 (n_213, in_0[6], in_1[3]);
  and g32 (n_247, in_0[7], in_1[3]);
  and g33 (n_63, in_0[0], in_1[4]);
  and g34 (n_83, in_0[1], in_1[4]);
  and g35 (n_109, in_0[2], in_1[4]);
  and g36 (n_142, in_0[3], in_1[4]);
  and g37 (n_176, in_0[4], in_1[4]);
  and g38 (n_220, in_0[5], in_1[4]);
  and g39 (n_248, in_0[6], in_1[4]);
  and g40 (n_277, in_0[7], in_1[4]);
  and g41 (n_87, in_0[0], in_1[5]);
  and g42 (n_113, in_0[1], in_1[5]);
  and g43 (n_146, in_0[2], in_1[5]);
  and g44 (n_179, in_0[3], in_1[5]);
  and g45 (n_214, in_0[4], in_1[5]);
  and g46 (n_254, in_0[5], in_1[5]);
  and g47 (n_278, in_0[6], in_1[5]);
  and g48 (n_301, in_0[7], in_1[5]);
  and g49 (n_116, in_0[0], in_1[6]);
  and g50 (n_149, in_0[1], in_1[6]);
  and g51 (n_183, in_0[2], in_1[6]);
  and g52 (n_217, in_0[3], in_1[6]);
  and g53 (n_249, in_0[4], in_1[6]);
  and g54 (n_282, in_0[5], in_1[6]);
  and g55 (n_302, in_0[6], in_1[6]);
  and g56 (n_319, in_0[7], in_1[6]);
  and g57 (n_139, in_0[0], in_1[7]);
  and g58 (n_186, in_0[1], in_1[7]);
  and g59 (n_221, in_0[2], in_1[7]);
  and g60 (n_252, in_0[3], in_1[7]);
  and g61 (n_279, in_0[4], in_1[7]);
  and g62 (n_305, in_0[5], in_1[7]);
  and g63 (n_320, in_0[6], in_1[7]);
  and g64 (n_331, in_0[7], in_1[7]);
  and g65 (out_1[0], in_2[0], in_3[0]);
  and g66 (n_35, in_2[1], in_3[0]);
  and g67 (n_39, in_2[2], in_3[0]);
  and g68 (n_48, in_2[3], in_3[0]);
  and g69 (n_66, in_2[4], in_3[0]);
  and g70 (n_89, in_2[5], in_3[0]);
  and g71 (n_107, in_2[6], in_3[0]);
  and g72 (n_141, in_2[7], in_3[0]);
  and g73 (n_34, in_2[0], in_3[1]);
  and g74 (n_40, in_2[1], in_3[1]);
  and g75 (n_50, in_2[2], in_3[1]);
  and g76 (n_67, in_2[3], in_3[1]);
  and g77 (n_81, in_2[4], in_3[1]);
  and g78 (n_108, in_2[5], in_3[1]);
  and g79 (n_143, in_2[6], in_3[1]);
  and g80 (n_177, in_2[7], in_3[1]);
  and g81 (n_38, in_2[0], in_3[2]);
  and g82 (n_51, in_2[1], in_3[2]);
  and g83 (n_61, in_2[2], in_3[2]);
  and g84 (n_82, in_2[3], in_3[2]);
  and g85 (n_110, in_2[4], in_3[2]);
  and g86 (n_144, in_2[5], in_3[2]);
  and g87 (n_178, in_2[6], in_3[2]);
  and g88 (n_223, in_2[7], in_3[2]);
  and g89 (n_47, in_2[0], in_3[3]);
  and g90 (n_62, in_2[1], in_3[3]);
  and g91 (n_84, in_2[2], in_3[3]);
  and g92 (n_111, in_2[3], in_3[3]);
  and g93 (n_147, in_2[4], in_3[3]);
  and g94 (n_180, in_2[5], in_3[3]);
  and g95 (n_215, in_2[6], in_3[3]);
  and g96 (n_255, in_2[7], in_3[3]);
  and g97 (n_64, in_2[0], in_3[4]);
  and g98 (n_85, in_2[1], in_3[4]);
  and g99 (n_114, in_2[2], in_3[4]);
  and g100 (n_148, in_2[3], in_3[4]);
  and g101 (n_181, in_2[4], in_3[4]);
  and g102 (n_216, in_2[5], in_3[4]);
  and g103 (n_256, in_2[6], in_3[4]);
  and g104 (n_281, in_2[7], in_3[4]);
  and g105 (n_88, in_2[0], in_3[5]);
  and g106 (n_115, in_2[1], in_3[5]);
  and g107 (n_150, in_2[2], in_3[5]);
  and g108 (n_184, in_2[3], in_3[5]);
  and g109 (n_218, in_2[4], in_3[5]);
  and g110 (n_250, in_2[5], in_3[5]);
  and g111 (n_283, in_2[6], in_3[5]);
  and g112 (n_303, in_2[7], in_3[5]);
  and g113 (n_117, in_2[0], in_3[6]);
  and g114 (n_151, in_2[1], in_3[6]);
  and g115 (n_185, in_2[2], in_3[6]);
  and g116 (n_219, in_2[3], in_3[6]);
  and g117 (n_251, in_2[4], in_3[6]);
  and g118 (n_284, in_2[5], in_3[6]);
  and g119 (n_304, in_2[6], in_3[6]);
  and g120 (n_322, in_2[7], in_3[6]);
  and g121 (n_140, in_2[0], in_3[7]);
  and g122 (n_187, in_2[1], in_3[7]);
  and g123 (n_222, in_2[2], in_3[7]);
  and g124 (n_253, in_2[3], in_3[7]);
  and g125 (n_280, in_2[4], in_3[7]);
  and g126 (n_306, in_2[5], in_3[7]);
  and g127 (n_321, in_2[6], in_3[7]);
  and g128 (n_332, in_2[7], in_3[7]);
  xor g233 (n_370, n_33, n_34);
  xor g234 (out_1[1], n_370, n_35);
  nand g235 (n_371, n_33, n_34);
  nand g236 (n_372, n_35, n_34);
  nand g237 (n_373, n_33, n_35);
  nand g238 (n_43, n_371, n_372, n_373);
  xor g239 (n_42, n_36, n_37);
  and g240 (n_52, n_36, n_37);
  xor g241 (n_374, n_38, n_39);
  xor g242 (out_0[2], n_374, n_40);
  nand g243 (n_375, n_38, n_39);
  nand g244 (n_376, n_40, n_39);
  nand g245 (n_377, n_38, n_40);
  nand g246 (n_54, n_375, n_376, n_377);
  xor g247 (n_378, n_41, n_42);
  xor g248 (out_1[2], n_378, n_43);
  nand g249 (n_379, n_41, n_42);
  nand g250 (n_380, n_43, n_42);
  nand g251 (n_381, n_41, n_43);
  nand g252 (out_0[3], n_379, n_380, n_381);
  xor g253 (n_53, n_44, n_45);
  and g254 (n_69, n_44, n_45);
  xor g255 (n_382, n_46, n_47);
  xor g256 (n_56, n_382, n_48);
  nand g257 (n_383, n_46, n_47);
  nand g258 (n_384, n_48, n_47);
  nand g259 (n_385, n_46, n_48);
  nand g260 (n_70, n_383, n_384, n_385);
  xor g261 (n_386, n_49, n_50);
  xor g262 (n_55, n_386, n_51);
  nand g263 (n_387, n_49, n_50);
  nand g264 (n_388, n_51, n_50);
  nand g265 (n_389, n_49, n_51);
  nand g266 (n_71, n_387, n_388, n_389);
  xor g267 (n_390, n_52, n_53);
  xor g268 (n_57, n_390, n_54);
  nand g269 (n_391, n_52, n_53);
  nand g270 (n_392, n_54, n_53);
  nand g271 (n_393, n_52, n_54);
  nand g272 (n_75, n_391, n_392, n_393);
  xor g273 (n_394, n_55, n_56);
  xor g274 (out_1[3], n_394, n_57);
  nand g275 (n_395, n_55, n_56);
  nand g276 (n_396, n_57, n_56);
  nand g277 (n_397, n_55, n_57);
  nand g278 (out_0[4], n_395, n_396, n_397);
  xor g279 (n_68, n_58, n_59);
  and g280 (n_91, n_58, n_59);
  xor g281 (n_398, n_60, n_61);
  xor g282 (n_72, n_398, n_62);
  nand g283 (n_399, n_60, n_61);
  nand g284 (n_400, n_62, n_61);
  nand g285 (n_401, n_60, n_62);
  nand g286 (n_93, n_399, n_400, n_401);
  xor g287 (n_402, n_63, n_64);
  xor g288 (n_73, n_402, n_65);
  nand g289 (n_403, n_63, n_64);
  nand g290 (n_404, n_65, n_64);
  nand g291 (n_405, n_63, n_65);
  nand g292 (n_92, n_403, n_404, n_405);
  xor g293 (n_406, n_66, n_67);
  xor g294 (n_74, n_406, n_68);
  nand g295 (n_407, n_66, n_67);
  nand g296 (n_408, n_68, n_67);
  nand g297 (n_409, n_66, n_68);
  nand g298 (n_97, n_407, n_408, n_409);
  xor g299 (n_410, n_69, n_70);
  xor g300 (n_76, n_410, n_71);
  nand g301 (n_411, n_69, n_70);
  nand g302 (n_412, n_71, n_70);
  nand g303 (n_413, n_69, n_71);
  nand g304 (n_98, n_411, n_412, n_413);
  xor g305 (n_414, n_72, n_73);
  xor g306 (n_77, n_414, n_74);
  nand g307 (n_415, n_72, n_73);
  nand g308 (n_416, n_74, n_73);
  nand g309 (n_417, n_72, n_74);
  nand g310 (n_101, n_415, n_416, n_417);
  xor g311 (n_418, n_75, n_76);
  xor g312 (out_1[4], n_418, n_77);
  nand g313 (n_419, n_75, n_76);
  nand g314 (n_420, n_77, n_76);
  nand g315 (n_421, n_75, n_77);
  nand g316 (out_0[5], n_419, n_420, n_421);
  xor g317 (n_90, n_78, n_79);
  and g318 (n_119, n_78, n_79);
  xor g319 (n_422, n_80, n_81);
  xor g320 (n_95, n_422, n_82);
  nand g321 (n_423, n_80, n_81);
  nand g322 (n_424, n_82, n_81);
  nand g323 (n_425, n_80, n_82);
  nand g324 (n_120, n_423, n_424, n_425);
  xor g325 (n_426, n_83, n_84);
  xor g326 (n_96, n_426, n_85);
  nand g327 (n_427, n_83, n_84);
  nand g328 (n_428, n_85, n_84);
  nand g329 (n_429, n_83, n_85);
  nand g330 (n_121, n_427, n_428, n_429);
  xor g331 (n_430, n_86, n_87);
  xor g332 (n_94, n_430, n_88);
  nand g333 (n_431, n_86, n_87);
  nand g334 (n_432, n_88, n_87);
  nand g335 (n_433, n_86, n_88);
  nand g336 (n_122, n_431, n_432, n_433);
  xor g337 (n_434, n_89, n_90);
  xor g338 (n_99, n_434, n_91);
  nand g339 (n_435, n_89, n_90);
  nand g340 (n_436, n_91, n_90);
  nand g341 (n_437, n_89, n_91);
  nand g342 (n_127, n_435, n_436, n_437);
  xor g343 (n_438, n_92, n_93);
  xor g344 (n_100, n_438, n_94);
  nand g345 (n_439, n_92, n_93);
  nand g346 (n_440, n_94, n_93);
  nand g347 (n_441, n_92, n_94);
  nand g348 (n_130, n_439, n_440, n_441);
  xor g349 (n_442, n_95, n_96);
  xor g350 (n_102, n_442, n_97);
  nand g351 (n_443, n_95, n_96);
  nand g352 (n_444, n_97, n_96);
  nand g353 (n_445, n_95, n_97);
  nand g354 (n_132, n_443, n_444, n_445);
  xor g355 (n_446, n_98, n_99);
  xor g356 (n_103, n_446, n_100);
  nand g357 (n_447, n_98, n_99);
  nand g358 (n_448, n_100, n_99);
  nand g359 (n_449, n_98, n_100);
  nand g360 (n_134, n_447, n_448, n_449);
  xor g361 (n_450, n_101, n_102);
  xor g362 (out_1[5], n_450, n_103);
  nand g363 (n_451, n_101, n_102);
  nand g364 (n_452, n_103, n_102);
  nand g365 (n_453, n_101, n_103);
  nand g366 (out_0[6], n_451, n_452, n_453);
  xor g367 (n_118, n_104, n_105);
  and g368 (n_152, n_104, n_105);
  xor g369 (n_454, n_106, n_107);
  xor g370 (n_123, n_454, n_108);
  nand g371 (n_455, n_106, n_107);
  nand g372 (n_456, n_108, n_107);
  nand g373 (n_457, n_106, n_108);
  nand g374 (n_154, n_455, n_456, n_457);
  xor g375 (n_458, n_109, n_110);
  xor g376 (n_125, n_458, n_111);
  nand g377 (n_459, n_109, n_110);
  nand g378 (n_460, n_111, n_110);
  nand g379 (n_461, n_109, n_111);
  nand g380 (n_157, n_459, n_460, n_461);
  xor g381 (n_462, n_112, n_113);
  xor g382 (n_126, n_462, n_114);
  nand g383 (n_463, n_112, n_113);
  nand g384 (n_464, n_114, n_113);
  nand g385 (n_465, n_112, n_114);
  nand g386 (n_155, n_463, n_464, n_465);
  xor g387 (n_466, n_115, n_116);
  xor g388 (n_124, n_466, n_117);
  nand g389 (n_467, n_115, n_116);
  nand g390 (n_468, n_117, n_116);
  nand g391 (n_469, n_115, n_117);
  nand g392 (n_156, n_467, n_468, n_469);
  xor g393 (n_470, n_118, n_119);
  xor g394 (n_128, n_470, n_120);
  nand g395 (n_471, n_118, n_119);
  nand g396 (n_472, n_120, n_119);
  nand g397 (n_473, n_118, n_120);
  nand g398 (n_163, n_471, n_472, n_473);
  xor g399 (n_474, n_121, n_122);
  xor g400 (n_129, n_474, n_123);
  nand g401 (n_475, n_121, n_122);
  nand g402 (n_476, n_123, n_122);
  nand g403 (n_477, n_121, n_123);
  nand g404 (n_165, n_475, n_476, n_477);
  xor g405 (n_478, n_124, n_125);
  xor g406 (n_131, n_478, n_126);
  nand g407 (n_479, n_124, n_125);
  nand g408 (n_480, n_126, n_125);
  nand g409 (n_481, n_124, n_126);
  nand g410 (n_164, n_479, n_480, n_481);
  xor g411 (n_482, n_127, n_128);
  xor g412 (n_133, n_482, n_129);
  nand g413 (n_483, n_127, n_128);
  nand g414 (n_484, n_129, n_128);
  nand g415 (n_485, n_127, n_129);
  nand g416 (n_169, n_483, n_484, n_485);
  xor g417 (n_486, n_130, n_131);
  xor g418 (n_135, n_486, n_132);
  nand g419 (n_487, n_130, n_131);
  nand g420 (n_488, n_132, n_131);
  nand g421 (n_489, n_130, n_132);
  nand g422 (n_172, n_487, n_488, n_489);
  xor g423 (n_490, n_133, n_134);
  xor g424 (out_1[6], n_490, n_135);
  nand g425 (n_491, n_133, n_134);
  nand g426 (n_492, n_135, n_134);
  nand g427 (n_493, n_133, n_135);
  nand g428 (out_0[7], n_491, n_492, n_493);
  xor g429 (n_153, n_136, n_137);
  and g430 (n_189, n_136, n_137);
  xor g431 (n_494, n_138, n_139);
  xor g432 (n_159, n_494, n_140);
  nand g433 (n_495, n_138, n_139);
  nand g434 (n_496, n_140, n_139);
  nand g435 (n_497, n_138, n_140);
  nand g436 (n_190, n_495, n_496, n_497);
  xor g437 (n_498, n_141, n_142);
  xor g438 (n_160, n_498, n_143);
  nand g439 (n_499, n_141, n_142);
  nand g440 (n_500, n_143, n_142);
  nand g441 (n_501, n_141, n_143);
  nand g442 (n_191, n_499, n_500, n_501);
  xor g443 (n_502, n_144, n_145);
  xor g444 (n_158, n_502, n_146);
  nand g445 (n_503, n_144, n_145);
  nand g446 (n_504, n_146, n_145);
  nand g447 (n_505, n_144, n_146);
  nand g448 (n_192, n_503, n_504, n_505);
  xor g449 (n_506, n_147, n_148);
  xor g450 (n_161, n_506, n_149);
  nand g451 (n_507, n_147, n_148);
  nand g452 (n_508, n_149, n_148);
  nand g453 (n_509, n_147, n_149);
  nand g454 (n_193, n_507, n_508, n_509);
  xor g455 (n_510, n_150, n_151);
  xor g456 (n_162, n_510, n_152);
  nand g457 (n_511, n_150, n_151);
  nand g458 (n_512, n_152, n_151);
  nand g459 (n_513, n_150, n_152);
  nand g460 (n_198, n_511, n_512, n_513);
  xor g461 (n_514, n_153, n_154);
  xor g462 (n_166, n_514, n_155);
  nand g463 (n_515, n_153, n_154);
  nand g464 (n_516, n_155, n_154);
  nand g465 (n_517, n_153, n_155);
  nand g466 (n_200, n_515, n_516, n_517);
  xor g467 (n_518, n_156, n_157);
  xor g468 (n_167, n_518, n_158);
  nand g469 (n_519, n_156, n_157);
  nand g470 (n_520, n_158, n_157);
  nand g471 (n_521, n_156, n_158);
  nand g472 (n_201, n_519, n_520, n_521);
  xor g473 (n_522, n_159, n_160);
  xor g474 (n_168, n_522, n_161);
  nand g475 (n_523, n_159, n_160);
  nand g476 (n_524, n_161, n_160);
  nand g477 (n_525, n_159, n_161);
  nand g478 (n_202, n_523, n_524, n_525);
  xor g479 (n_526, n_162, n_163);
  xor g480 (n_170, n_526, n_164);
  nand g481 (n_527, n_162, n_163);
  nand g482 (n_528, n_164, n_163);
  nand g483 (n_529, n_162, n_164);
  nand g484 (n_207, n_527, n_528, n_529);
  xor g485 (n_530, n_165, n_166);
  xor g486 (n_171, n_530, n_167);
  nand g487 (n_531, n_165, n_166);
  nand g488 (n_532, n_167, n_166);
  nand g489 (n_533, n_165, n_167);
  nand g490 (n_206, n_531, n_532, n_533);
  xor g491 (n_534, n_168, n_169);
  xor g492 (n_173, n_534, n_170);
  nand g493 (n_535, n_168, n_169);
  nand g494 (n_536, n_170, n_169);
  nand g495 (n_537, n_168, n_170);
  nand g496 (n_210, n_535, n_536, n_537);
  xor g497 (n_538, n_171, n_172);
  xor g498 (out_1[7], n_538, n_173);
  nand g499 (n_539, n_171, n_172);
  nand g500 (n_540, n_173, n_172);
  nand g501 (n_541, n_171, n_173);
  nand g502 (out_0[8], n_539, n_540, n_541);
  xor g503 (n_188, n_174, n_175);
  and g504 (n_225, n_174, n_175);
  xor g505 (n_542, n_176, n_177);
  xor g506 (n_194, n_542, n_178);
  nand g507 (n_543, n_176, n_177);
  nand g508 (n_544, n_178, n_177);
  nand g509 (n_545, n_176, n_178);
  nand g510 (n_228, n_543, n_544, n_545);
  xor g511 (n_546, n_179, n_180);
  xor g512 (n_196, n_546, n_181);
  nand g513 (n_547, n_179, n_180);
  nand g514 (n_548, n_181, n_180);
  nand g515 (n_549, n_179, n_181);
  nand g516 (n_229, n_547, n_548, n_549);
  xor g517 (n_550, n_182, n_183);
  xor g518 (n_195, n_550, n_184);
  nand g519 (n_551, n_182, n_183);
  nand g520 (n_552, n_184, n_183);
  nand g521 (n_553, n_182, n_184);
  nand g522 (n_226, n_551, n_552, n_553);
  xor g523 (n_554, n_185, n_186);
  xor g524 (n_197, n_554, n_187);
  nand g525 (n_555, n_185, n_186);
  nand g526 (n_556, n_187, n_186);
  nand g527 (n_557, n_185, n_187);
  nand g528 (n_227, n_555, n_556, n_557);
  xor g529 (n_558, n_188, n_189);
  xor g530 (n_199, n_558, n_190);
  nand g531 (n_559, n_188, n_189);
  nand g532 (n_560, n_190, n_189);
  nand g533 (n_561, n_188, n_190);
  nand g534 (n_234, n_559, n_560, n_561);
  xor g535 (n_562, n_191, n_192);
  xor g536 (n_203, n_562, n_193);
  nand g537 (n_563, n_191, n_192);
  nand g538 (n_564, n_193, n_192);
  nand g539 (n_565, n_191, n_193);
  nand g540 (n_235, n_563, n_564, n_565);
  xor g541 (n_566, n_194, n_195);
  xor g542 (n_204, n_566, n_196);
  nand g543 (n_567, n_194, n_195);
  nand g544 (n_568, n_196, n_195);
  nand g545 (n_569, n_194, n_196);
  nand g546 (n_236, n_567, n_568, n_569);
  xor g547 (n_570, n_197, n_198);
  xor g548 (n_205, n_570, n_199);
  nand g549 (n_571, n_197, n_198);
  nand g550 (n_572, n_199, n_198);
  nand g551 (n_573, n_197, n_199);
  nand g552 (n_239, n_571, n_572, n_573);
  xor g553 (n_574, n_200, n_201);
  xor g554 (n_208, n_574, n_202);
  nand g555 (n_575, n_200, n_201);
  nand g556 (n_576, n_202, n_201);
  nand g557 (n_577, n_200, n_202);
  nand g558 (n_240, n_575, n_576, n_577);
  xor g559 (n_578, n_203, n_204);
  xor g560 (n_209, n_578, n_205);
  nand g561 (n_579, n_203, n_204);
  nand g562 (n_580, n_205, n_204);
  nand g563 (n_581, n_203, n_205);
  nand g564 (n_243, n_579, n_580, n_581);
  xor g565 (n_582, n_206, n_207);
  xor g566 (n_211, n_582, n_208);
  nand g567 (n_583, n_206, n_207);
  nand g568 (n_584, n_208, n_207);
  nand g569 (n_585, n_206, n_208);
  nand g570 (n_245, n_583, n_584, n_585);
  xor g571 (n_586, n_209, n_210);
  xor g572 (out_1[8], n_586, n_211);
  nand g573 (n_587, n_209, n_210);
  nand g574 (n_588, n_211, n_210);
  nand g575 (n_589, n_209, n_211);
  nand g576 (out_0[9], n_587, n_588, n_589);
  xor g577 (n_224, n_212, n_213);
  and g578 (n_257, n_212, n_213);
  xor g579 (n_590, n_214, n_215);
  xor g580 (n_231, n_590, n_216);
  nand g581 (n_591, n_214, n_215);
  nand g582 (n_592, n_216, n_215);
  nand g583 (n_593, n_214, n_216);
  nand g584 (n_258, n_591, n_592, n_593);
  xor g585 (n_594, n_217, n_218);
  xor g586 (n_232, n_594, n_219);
  nand g587 (n_595, n_217, n_218);
  nand g588 (n_596, n_219, n_218);
  nand g589 (n_597, n_217, n_219);
  nand g590 (n_259, n_595, n_596, n_597);
  xor g591 (n_598, n_220, n_221);
  xor g592 (n_230, n_598, n_222);
  nand g593 (n_599, n_220, n_221);
  nand g594 (n_600, n_222, n_221);
  nand g595 (n_601, n_220, n_222);
  nand g596 (n_260, n_599, n_600, n_601);
  xor g597 (n_602, n_223, n_224);
  xor g598 (n_233, n_602, n_225);
  nand g599 (n_603, n_223, n_224);
  nand g600 (n_604, n_225, n_224);
  nand g601 (n_605, n_223, n_225);
  nand g602 (n_264, n_603, n_604, n_605);
  xor g603 (n_606, n_226, n_227);
  xor g604 (n_237, n_606, n_228);
  nand g605 (n_607, n_226, n_227);
  nand g606 (n_608, n_228, n_227);
  nand g607 (n_609, n_226, n_228);
  nand g608 (n_265, n_607, n_608, n_609);
  xor g609 (n_610, n_229, n_230);
  xor g610 (n_238, n_610, n_231);
  nand g611 (n_611, n_229, n_230);
  nand g612 (n_612, n_231, n_230);
  nand g613 (n_613, n_229, n_231);
  nand g614 (n_267, n_611, n_612, n_613);
  xor g615 (n_614, n_232, n_233);
  xor g616 (n_241, n_614, n_234);
  nand g617 (n_615, n_232, n_233);
  nand g618 (n_616, n_234, n_233);
  nand g619 (n_617, n_232, n_234);
  nand g620 (n_270, n_615, n_616, n_617);
  xor g621 (n_618, n_235, n_236);
  xor g622 (n_242, n_618, n_237);
  nand g623 (n_619, n_235, n_236);
  nand g624 (n_620, n_237, n_236);
  nand g625 (n_621, n_235, n_237);
  nand g626 (n_272, n_619, n_620, n_621);
  xor g627 (n_622, n_238, n_239);
  xor g628 (n_244, n_622, n_240);
  nand g629 (n_623, n_238, n_239);
  nand g630 (n_624, n_240, n_239);
  nand g631 (n_625, n_238, n_240);
  nand g632 (n_274, n_623, n_624, n_625);
  xor g633 (n_626, n_241, n_242);
  xor g634 (n_246, n_626, n_243);
  nand g635 (n_627, n_241, n_242);
  nand g636 (n_628, n_243, n_242);
  nand g637 (n_629, n_241, n_243);
  nand g638 (n_276, n_627, n_628, n_629);
  xor g639 (n_630, n_244, n_245);
  xor g640 (out_1[9], n_630, n_246);
  nand g641 (n_631, n_244, n_245);
  nand g642 (n_632, n_246, n_245);
  nand g643 (n_633, n_244, n_246);
  nand g644 (out_0[10], n_631, n_632, n_633);
  xor g645 (n_634, n_247, n_248);
  xor g646 (n_263, n_634, n_249);
  nand g647 (n_635, n_247, n_248);
  nand g648 (n_636, n_249, n_248);
  nand g649 (n_637, n_247, n_249);
  nand g650 (n_285, n_635, n_636, n_637);
  xor g651 (n_638, n_250, n_251);
  xor g652 (n_261, n_638, n_252);
  nand g653 (n_639, n_250, n_251);
  nand g654 (n_640, n_252, n_251);
  nand g655 (n_641, n_250, n_252);
  nand g656 (n_286, n_639, n_640, n_641);
  xor g657 (n_642, n_253, n_254);
  xor g658 (n_262, n_642, n_255);
  nand g659 (n_643, n_253, n_254);
  nand g660 (n_644, n_255, n_254);
  nand g661 (n_645, n_253, n_255);
  nand g662 (n_287, n_643, n_644, n_645);
  xor g663 (n_646, n_256, n_257);
  xor g664 (n_266, n_646, n_258);
  nand g665 (n_647, n_256, n_257);
  nand g666 (n_648, n_258, n_257);
  nand g667 (n_649, n_256, n_258);
  nand g668 (n_291, n_647, n_648, n_649);
  xor g669 (n_650, n_259, n_260);
  xor g670 (n_268, n_650, n_261);
  nand g671 (n_651, n_259, n_260);
  nand g672 (n_652, n_261, n_260);
  nand g673 (n_653, n_259, n_261);
  nand g674 (n_293, n_651, n_652, n_653);
  xor g675 (n_654, n_262, n_263);
  xor g676 (n_269, n_654, n_264);
  nand g677 (n_655, n_262, n_263);
  nand g678 (n_656, n_264, n_263);
  nand g679 (n_657, n_262, n_264);
  nand g680 (n_294, n_655, n_656, n_657);
  xor g681 (n_658, n_265, n_266);
  xor g682 (n_271, n_658, n_267);
  nand g683 (n_659, n_265, n_266);
  nand g684 (n_660, n_267, n_266);
  nand g685 (n_661, n_265, n_267);
  nand g686 (n_296, n_659, n_660, n_661);
  xor g687 (n_662, n_268, n_269);
  xor g688 (n_273, n_662, n_270);
  nand g689 (n_663, n_268, n_269);
  nand g690 (n_664, n_270, n_269);
  nand g691 (n_665, n_268, n_270);
  nand g692 (n_298, n_663, n_664, n_665);
  xor g693 (n_666, n_271, n_272);
  xor g694 (n_275, n_666, n_273);
  nand g695 (n_667, n_271, n_272);
  nand g696 (n_668, n_273, n_272);
  nand g697 (n_669, n_271, n_273);
  nand g698 (n_300, n_667, n_668, n_669);
  xor g699 (n_670, n_274, n_275);
  xor g700 (out_1[10], n_670, n_276);
  nand g701 (n_671, n_274, n_275);
  nand g702 (n_672, n_276, n_275);
  nand g703 (n_673, n_274, n_276);
  nand g704 (out_0[11], n_671, n_672, n_673);
  xor g705 (n_674, n_277, n_278);
  xor g706 (n_288, n_674, n_279);
  nand g707 (n_675, n_277, n_278);
  nand g708 (n_676, n_279, n_278);
  nand g709 (n_677, n_277, n_279);
  nand g710 (n_308, n_675, n_676, n_677);
  xor g711 (n_678, n_280, n_281);
  xor g712 (n_289, n_678, n_282);
  nand g713 (n_679, n_280, n_281);
  nand g714 (n_680, n_282, n_281);
  nand g715 (n_681, n_280, n_282);
  nand g716 (n_307, n_679, n_680, n_681);
  xor g717 (n_682, n_283, n_284);
  xor g718 (n_290, n_682, n_285);
  nand g719 (n_683, n_283, n_284);
  nand g720 (n_684, n_285, n_284);
  nand g721 (n_685, n_283, n_285);
  nand g722 (n_311, n_683, n_684, n_685);
  xor g723 (n_686, n_286, n_287);
  xor g724 (n_292, n_686, n_288);
  nand g725 (n_687, n_286, n_287);
  nand g726 (n_688, n_288, n_287);
  nand g727 (n_689, n_286, n_288);
  nand g728 (n_313, n_687, n_688, n_689);
  xor g729 (n_690, n_289, n_290);
  xor g730 (n_295, n_690, n_291);
  nand g731 (n_691, n_289, n_290);
  nand g732 (n_692, n_291, n_290);
  nand g733 (n_693, n_289, n_291);
  nand g734 (n_314, n_691, n_692, n_693);
  xor g735 (n_694, n_292, n_293);
  xor g736 (n_297, n_694, n_294);
  nand g737 (n_695, n_292, n_293);
  nand g738 (n_696, n_294, n_293);
  nand g739 (n_697, n_292, n_294);
  nand g740 (n_316, n_695, n_696, n_697);
  xor g741 (n_698, n_295, n_296);
  xor g742 (n_299, n_698, n_297);
  nand g743 (n_699, n_295, n_296);
  nand g744 (n_700, n_297, n_296);
  nand g745 (n_701, n_295, n_297);
  nand g746 (n_318, n_699, n_700, n_701);
  xor g747 (n_702, n_298, n_299);
  xor g748 (out_1[11], n_702, n_300);
  nand g749 (n_703, n_298, n_299);
  nand g750 (n_704, n_300, n_299);
  nand g751 (n_705, n_298, n_300);
  nand g752 (out_1[12], n_703, n_704, n_705);
  xor g753 (n_706, n_301, n_302);
  xor g754 (n_310, n_706, n_303);
  nand g755 (n_707, n_301, n_302);
  nand g756 (n_708, n_303, n_302);
  nand g757 (n_709, n_301, n_303);
  nand g758 (n_323, n_707, n_708, n_709);
  xor g759 (n_710, n_304, n_305);
  xor g760 (n_309, n_710, n_306);
  nand g761 (n_711, n_304, n_305);
  nand g762 (n_712, n_306, n_305);
  nand g763 (n_713, n_304, n_306);
  nand g764 (n_324, n_711, n_712, n_713);
  xor g765 (n_714, n_307, n_308);
  xor g766 (n_312, n_714, n_309);
  nand g767 (n_715, n_307, n_308);
  nand g768 (n_716, n_309, n_308);
  nand g769 (n_717, n_307, n_309);
  nand g770 (n_327, n_715, n_716, n_717);
  xor g771 (n_718, n_310, n_311);
  xor g772 (n_315, n_718, n_312);
  nand g773 (n_719, n_310, n_311);
  nand g774 (n_720, n_312, n_311);
  nand g775 (n_721, n_310, n_312);
  nand g776 (n_328, n_719, n_720, n_721);
  xor g777 (n_722, n_313, n_314);
  xor g778 (n_317, n_722, n_315);
  nand g779 (n_723, n_313, n_314);
  nand g780 (n_724, n_315, n_314);
  nand g781 (n_725, n_313, n_315);
  nand g782 (n_330, n_723, n_724, n_725);
  xor g783 (n_726, n_316, n_317);
  xor g784 (out_0[12], n_726, n_318);
  nand g785 (n_727, n_316, n_317);
  nand g786 (n_728, n_318, n_317);
  nand g787 (n_729, n_316, n_318);
  nand g788 (out_1[13], n_727, n_728, n_729);
  xor g789 (n_730, n_319, n_320);
  xor g790 (n_325, n_730, n_321);
  nand g791 (n_731, n_319, n_320);
  nand g792 (n_732, n_321, n_320);
  nand g793 (n_733, n_319, n_321);
  nand g794 (n_333, n_731, n_732, n_733);
  xor g795 (n_734, n_322, n_323);
  xor g796 (n_326, n_734, n_324);
  nand g797 (n_735, n_322, n_323);
  nand g798 (n_736, n_324, n_323);
  nand g799 (n_737, n_322, n_324);
  nand g800 (n_334, n_735, n_736, n_737);
  xor g801 (n_738, n_325, n_326);
  xor g802 (n_329, n_738, n_327);
  nand g803 (n_739, n_325, n_326);
  nand g804 (n_740, n_327, n_326);
  nand g805 (n_741, n_325, n_327);
  nand g806 (n_336, n_739, n_740, n_741);
  xor g807 (n_742, n_328, n_329);
  xor g808 (out_0[13], n_742, n_330);
  nand g809 (n_743, n_328, n_329);
  nand g810 (n_744, n_330, n_329);
  nand g811 (n_745, n_328, n_330);
  nand g812 (out_1[14], n_743, n_744, n_745);
  xor g813 (n_746, n_331, n_332);
  xor g814 (n_335, n_746, n_333);
  nand g815 (n_747, n_331, n_332);
  nand g816 (n_748, n_333, n_332);
  nand g817 (n_749, n_331, n_333);
  nand g818 (out_0[15], n_747, n_748, n_749);
  xor g819 (n_750, n_334, n_335);
  xor g820 (out_0[14], n_750, n_336);
  nand g821 (n_751, n_334, n_335);
  nand g822 (n_752, n_336, n_335);
  nand g823 (n_753, n_334, n_336);
  nand g824 (out_1[15], n_751, n_752, n_753);
endmodule

module csa_tree_GENERIC(in_0, in_1, in_2, in_3, out_0, out_1);
  input [7:0] in_0, in_1, in_2, in_3;
  output [16:0] out_0, out_1;
  wire [7:0] in_0, in_1, in_2, in_3;
  wire [16:0] out_0, out_1;
  csa_tree_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2 (in_2),
       .in_3 (in_3), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_add_25_30_group_50_GENERIC_REAL(in_0, in_1, in_2, in_3,
     out_0);
// synthesis_equation "assign out_0 = ( ( in_2 + in_3 ) + ( in_0 * in_1 )  )  ;"
  input [16:0] in_0, in_2, in_3;
  input [7:0] in_1;
  output [16:0] out_0;
  wire [16:0] in_0, in_2, in_3;
  wire [7:0] in_1;
  wire [16:0] out_0;
  wire n_43, n_60, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_115, n_116, n_117;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_172, n_174;
  wire n_175, n_176, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_221, n_223, n_224, n_225, n_227, n_228;
  wire n_229, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_270, n_272, n_273;
  wire n_274, n_276, n_277, n_278, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_313, n_315, n_316, n_326, n_329, n_332;
  wire n_335, n_338, n_341, n_344, n_347, n_354, n_355, n_356;
  wire n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364;
  wire n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372;
  wire n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380;
  wire n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_416, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_456, n_457, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_498, n_499;
  wire n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_510, n_511, n_512, n_513, n_514, n_515, n_516;
  wire n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532;
  wire n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540;
  wire n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548;
  wire n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556;
  wire n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564;
  wire n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572;
  wire n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580;
  wire n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588;
  wire n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596;
  wire n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604;
  wire n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_614;
  wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_640;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_660, n_662, n_663, n_664, n_665, n_666, n_667, n_668;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_680, n_682, n_683, n_684, n_685, n_686, n_687;
  wire n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695;
  wire n_696, n_697, n_700, n_702, n_703, n_704, n_705, n_706;
  wire n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714;
  wire n_715, n_716, n_717, n_720, n_722, n_723, n_724, n_725;
  wire n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733;
  wire n_734, n_735, n_736, n_737, n_740, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_758, n_762;
  wire n_766, n_767, n_768, n_769, n_770, n_772, n_774, n_775;
  wire n_777, n_779, n_780, n_782, n_784, n_785, n_787, n_789;
  wire n_790, n_792, n_794, n_795, n_797, n_799, n_800, n_802;
  wire n_804, n_805, n_807, n_809, n_810, n_812, n_814, n_815;
  wire n_817, n_819, n_820, n_822, n_824, n_825, n_827, n_829;
  wire n_830, n_832, n_834, n_835, n_837, n_839, n_840, n_842;
  wire n_844, n_845, n_847, n_864, n_867, n_868, n_869, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924;
  xor g2 (n_115, in_1[1], in_1[0]);
  xor g8 (n_116, in_1[1], in_0[0]);
  and g12 (n_110, in_0[0], in_1[0]);
  xor g13 (n_121, in_1[1], in_0[1]);
  nand g14 (n_122, n_121, in_1[0]);
  nand g15 (n_123, n_116, n_117);
  nand g16 (n_92, n_122, n_123);
  xor g17 (n_124, in_1[1], in_0[2]);
  nand g18 (n_125, n_124, in_1[0]);
  nand g19 (n_126, n_121, n_117);
  nand g20 (n_357, n_125, n_126);
  xor g21 (n_127, in_1[1], in_0[3]);
  nand g22 (n_128, n_127, in_1[0]);
  nand g23 (n_129, n_124, n_117);
  nand g24 (n_361, n_128, n_129);
  xor g25 (n_130, in_1[1], in_0[4]);
  nand g26 (n_131, n_130, in_1[0]);
  nand g27 (n_132, n_127, n_117);
  nand g28 (n_368, n_131, n_132);
  xor g29 (n_133, in_1[1], in_0[5]);
  nand g30 (n_134, n_133, in_1[0]);
  nand g31 (n_135, n_130, n_117);
  nand g32 (n_373, n_134, n_135);
  xor g33 (n_136, in_1[1], in_0[6]);
  nand g34 (n_137, n_136, in_1[0]);
  nand g35 (n_138, n_133, n_117);
  nand g36 (n_383, n_137, n_138);
  xor g37 (n_139, in_1[1], in_0[7]);
  nand g38 (n_140, n_139, in_1[0]);
  nand g39 (n_141, n_136, n_117);
  nand g40 (n_396, n_140, n_141);
  xor g41 (n_142, in_1[1], in_0[8]);
  nand g42 (n_43, n_142, in_1[0]);
  nand g43 (n_143, n_139, n_117);
  nand g44 (n_408, n_43, n_143);
  xor g45 (n_144, in_1[1], in_0[9]);
  nand g46 (n_145, n_144, in_1[0]);
  nand g47 (n_146, n_142, n_117);
  nand g48 (n_420, n_145, n_146);
  xor g49 (n_147, in_1[1], in_0[10]);
  nand g50 (n_148, n_147, in_1[0]);
  nand g51 (n_149, n_144, n_117);
  nand g52 (n_431, n_148, n_149);
  xor g53 (n_150, in_1[1], in_0[11]);
  nand g54 (n_151, n_150, in_1[0]);
  nand g55 (n_152, n_147, n_117);
  nand g56 (n_444, n_151, n_152);
  xor g57 (n_153, in_1[1], in_0[12]);
  nand g58 (n_154, n_153, in_1[0]);
  nand g59 (n_60, n_150, n_117);
  nand g60 (n_457, n_154, n_60);
  xor g61 (n_155, in_1[1], in_0[13]);
  nand g62 (n_156, n_155, in_1[0]);
  nand g63 (n_157, n_153, n_117);
  nand g64 (n_470, n_156, n_157);
  xor g65 (n_158, in_1[1], in_0[14]);
  nand g66 (n_159, n_158, in_1[0]);
  nand g67 (n_160, n_155, n_117);
  nand g68 (n_483, n_159, n_160);
  xor g69 (n_161, in_1[1], in_0[15]);
  nand g70 (n_162, n_161, in_1[0]);
  nand g71 (n_163, n_158, n_117);
  nand g72 (n_496, n_162, n_163);
  xor g73 (n_164, in_1[1], in_0[16]);
  nand g74 (n_165, n_164, in_1[0]);
  nand g75 (n_166, n_161, n_117);
  nand g76 (n_508, n_165, n_166);
  xor g81 (n_172, in_1[2], in_1[1]);
  xor g82 (n_174, in_1[3], in_1[2]);
  nor g86 (n_223, in_1[1], in_1[2]);
  nand g87 (n_221, in_1[1], in_1[2]);
  xor g88 (n_175, in_1[3], in_0[0]);
  and g92 (n_356, in_0[0], n_172);
  xor g93 (n_180, in_1[3], in_0[1]);
  nand g94 (n_93, n_180, n_172);
  nand g95 (n_181, n_175, n_176);
  nand g96 (n_362, n_93, n_181);
  xor g97 (n_182, in_1[3], in_0[2]);
  nand g98 (n_183, n_182, n_172);
  nand g99 (n_184, n_180, n_176);
  nand g100 (n_367, n_183, n_184);
  xor g101 (n_185, in_1[3], in_0[3]);
  nand g102 (n_186, n_185, n_172);
  nand g103 (n_187, n_182, n_176);
  nand g104 (n_375, n_186, n_187);
  xor g105 (n_188, in_1[3], in_0[4]);
  nand g106 (n_189, n_188, n_172);
  nand g107 (n_190, n_185, n_176);
  nand g108 (n_382, n_189, n_190);
  xor g109 (n_191, in_1[3], in_0[5]);
  nand g110 (n_192, n_191, n_172);
  nand g111 (n_193, n_188, n_176);
  nand g112 (n_395, n_192, n_193);
  xor g113 (n_194, in_1[3], in_0[6]);
  nand g114 (n_195, n_194, n_172);
  nand g115 (n_196, n_191, n_176);
  nand g116 (n_407, n_195, n_196);
  xor g117 (n_197, in_1[3], in_0[7]);
  nand g118 (n_111, n_197, n_172);
  nand g119 (n_198, n_194, n_176);
  nand g120 (n_416, n_111, n_198);
  xor g121 (n_199, in_1[3], in_0[8]);
  nand g122 (n_200, n_199, n_172);
  nand g123 (n_201, n_197, n_176);
  nand g124 (n_428, n_200, n_201);
  xor g125 (n_202, in_1[3], in_0[9]);
  nand g126 (n_203, n_202, n_172);
  nand g127 (n_204, n_199, n_176);
  nand g128 (n_441, n_203, n_204);
  xor g129 (n_205, in_1[3], in_0[10]);
  nand g130 (n_206, n_205, n_172);
  nand g131 (n_207, n_202, n_176);
  nand g132 (n_454, n_206, n_207);
  xor g133 (n_208, in_1[3], in_0[11]);
  nand g134 (n_209, n_208, n_172);
  nand g135 (n_210, n_205, n_176);
  nand g136 (n_467, n_209, n_210);
  xor g137 (n_211, in_1[3], in_0[12]);
  nand g138 (n_212, n_211, n_172);
  nand g139 (n_213, n_208, n_176);
  nand g140 (n_480, n_212, n_213);
  xor g141 (n_214, in_1[3], in_0[13]);
  nand g142 (n_215, n_214, n_172);
  nand g143 (n_216, n_211, n_176);
  nand g144 (n_493, n_215, n_216);
  xor g145 (n_217, in_1[3], in_0[14]);
  nand g146 (n_218, n_217, n_172);
  nand g147 (n_219, n_214, n_176);
  nand g148 (n_507, n_218, n_219);
  or g151 (n_224, n_867, n_223);
  and g152 (n_360, in_1[3], n_224);
  xor g153 (n_225, in_1[4], in_1[3]);
  xor g154 (n_227, in_1[5], in_1[4]);
  nor g158 (n_272, in_1[3], in_1[4]);
  nand g159 (n_270, in_1[3], in_1[4]);
  xor g160 (n_228, in_1[5], in_0[0]);
  and g164 (n_365, in_0[0], n_225);
  xor g165 (n_233, in_1[5], in_0[1]);
  nand g166 (n_234, n_233, n_225);
  nand g167 (n_235, n_228, n_229);
  nand g168 (n_376, n_234, n_235);
  xor g169 (n_236, in_1[5], in_0[2]);
  nand g170 (n_237, n_236, n_225);
  nand g171 (n_238, n_233, n_229);
  nand g172 (n_385, n_237, n_238);
  xor g173 (n_239, in_1[5], in_0[3]);
  nand g174 (n_240, n_239, n_225);
  nand g175 (n_241, n_236, n_229);
  nand g176 (n_394, n_240, n_241);
  xor g177 (n_242, in_1[5], in_0[4]);
  nand g178 (n_243, n_242, n_225);
  nand g179 (n_244, n_239, n_229);
  nand g180 (n_406, n_243, n_244);
  xor g181 (n_245, in_1[5], in_0[5]);
  nand g182 (n_246, n_245, n_225);
  nand g183 (n_247, n_242, n_229);
  nand g184 (n_419, n_246, n_247);
  xor g185 (n_248, in_1[5], in_0[6]);
  nand g186 (n_249, n_248, n_225);
  nand g187 (n_250, n_245, n_229);
  nand g188 (n_430, n_249, n_250);
  xor g189 (n_251, in_1[5], in_0[7]);
  nand g190 (n_252, n_251, n_225);
  nand g191 (n_253, n_248, n_229);
  nand g192 (n_443, n_252, n_253);
  xor g193 (n_254, in_1[5], in_0[8]);
  nand g194 (n_255, n_254, n_225);
  nand g195 (n_256, n_251, n_229);
  nand g196 (n_456, n_255, n_256);
  xor g197 (n_257, in_1[5], in_0[9]);
  nand g198 (n_258, n_257, n_225);
  nand g199 (n_259, n_254, n_229);
  nand g200 (n_469, n_258, n_259);
  xor g201 (n_260, in_1[5], in_0[10]);
  nand g202 (n_261, n_260, n_225);
  nand g203 (n_262, n_257, n_229);
  nand g204 (n_482, n_261, n_262);
  xor g205 (n_263, in_1[5], in_0[11]);
  nand g206 (n_264, n_263, n_225);
  nand g207 (n_265, n_260, n_229);
  nand g208 (n_495, n_264, n_265);
  xor g209 (n_266, in_1[5], in_0[12]);
  nand g210 (n_267, n_266, n_225);
  nand g211 (n_268, n_263, n_229);
  nand g212 (n_506, n_267, n_268);
  or g215 (n_273, n_868, n_272);
  and g216 (n_372, in_1[5], n_273);
  xor g217 (n_274, in_1[6], in_1[5]);
  xor g218 (n_276, in_1[7], in_1[6]);
  nor g222 (n_315, in_1[5], in_1[6]);
  nand g223 (n_313, in_1[5], in_1[6]);
  xor g224 (n_277, in_1[7], in_0[0]);
  and g228 (n_381, in_0[0], n_274);
  xor g229 (n_282, in_1[7], in_0[1]);
  nand g230 (n_283, n_282, n_274);
  nand g231 (n_284, n_277, n_278);
  nand g232 (n_393, n_283, n_284);
  xor g233 (n_285, in_1[7], in_0[2]);
  nand g234 (n_286, n_285, n_274);
  nand g235 (n_287, n_282, n_278);
  nand g236 (n_405, n_286, n_287);
  xor g237 (n_288, in_1[7], in_0[3]);
  nand g238 (n_289, n_288, n_274);
  nand g239 (n_290, n_285, n_278);
  nand g240 (n_418, n_289, n_290);
  xor g241 (n_291, in_1[7], in_0[4]);
  nand g242 (n_292, n_291, n_274);
  nand g243 (n_293, n_288, n_278);
  nand g244 (n_429, n_292, n_293);
  xor g245 (n_294, in_1[7], in_0[5]);
  nand g246 (n_295, n_294, n_274);
  nand g247 (n_296, n_291, n_278);
  nand g248 (n_442, n_295, n_296);
  xor g249 (n_297, in_1[7], in_0[6]);
  nand g250 (n_298, n_297, n_274);
  nand g251 (n_299, n_294, n_278);
  nand g252 (n_455, n_298, n_299);
  xor g253 (n_300, in_1[7], in_0[7]);
  nand g254 (n_301, n_300, n_274);
  nand g255 (n_302, n_297, n_278);
  nand g256 (n_468, n_301, n_302);
  xor g257 (n_303, in_1[7], in_0[8]);
  nand g258 (n_304, n_303, n_274);
  nand g259 (n_305, n_300, n_278);
  nand g260 (n_481, n_304, n_305);
  xor g261 (n_306, in_1[7], in_0[9]);
  nand g262 (n_307, n_306, n_274);
  nand g263 (n_308, n_303, n_278);
  nand g264 (n_494, n_307, n_308);
  xor g265 (n_309, in_1[7], in_0[10]);
  nand g266 (n_310, n_309, n_274);
  nand g267 (n_311, n_306, n_278);
  nand g268 (n_510, n_310, n_311);
  or g271 (n_316, n_869, n_315);
  and g272 (n_391, in_1[7], n_316);
  and g284 (n_403, in_0[0], in_1[7]);
  nand g286 (n_326, in_0[1], in_1[7]);
  nand g290 (n_329, in_0[2], in_1[7]);
  nand g294 (n_332, in_0[3], in_1[7]);
  nand g298 (n_335, in_0[4], in_1[7]);
  nand g302 (n_338, in_0[5], in_1[7]);
  nand g306 (n_341, in_0[6], in_1[7]);
  nand g310 (n_344, in_0[7], in_1[7]);
  nand g314 (n_347, in_0[8], in_1[7]);
  xor g387 (n_518, in_2[1], in_3[1]);
  xor g388 (n_109, n_518, n_354);
  nand g389 (n_519, in_2[1], in_3[1]);
  nand g390 (n_520, n_354, in_3[1]);
  nand g391 (n_521, in_2[1], n_354);
  nand g392 (n_91, n_519, n_520, n_521);
  xor g393 (n_355, in_2[2], in_3[2]);
  and g394 (n_358, in_2[2], in_3[2]);
  xor g395 (n_522, n_355, n_356);
  xor g396 (n_108, n_522, n_357);
  nand g397 (n_523, n_355, n_356);
  nand g398 (n_524, n_357, n_356);
  nand g399 (n_525, n_355, n_357);
  nand g400 (n_90, n_523, n_524, n_525);
  xor g401 (n_359, in_2[3], in_3[3]);
  and g402 (n_364, in_2[3], in_3[3]);
  xor g403 (n_526, n_358, n_359);
  xor g404 (n_363, n_526, n_360);
  nand g405 (n_527, n_358, n_359);
  nand g406 (n_528, n_360, n_359);
  nand g407 (n_529, n_358, n_360);
  nand g408 (n_369, n_527, n_528, n_529);
  xor g409 (n_530, n_361, n_362);
  xor g410 (n_107, n_530, n_363);
  nand g411 (n_531, n_361, n_362);
  nand g412 (n_532, n_363, n_362);
  nand g413 (n_533, n_361, n_363);
  nand g414 (n_370, n_531, n_532, n_533);
  xor g415 (n_534, in_2[4], in_3[4]);
  xor g416 (n_366, n_534, n_364);
  nand g417 (n_535, in_2[4], in_3[4]);
  nand g418 (n_536, n_364, in_3[4]);
  nand g419 (n_537, in_2[4], n_364);
  nand g420 (n_374, n_535, n_536, n_537);
  xor g421 (n_538, n_365, n_366);
  xor g422 (n_89, n_538, n_367);
  nand g423 (n_539, n_365, n_366);
  nand g424 (n_540, n_367, n_366);
  nand g425 (n_541, n_365, n_367);
  nand g426 (n_377, n_539, n_540, n_541);
  xor g427 (n_542, n_368, n_369);
  xor g428 (n_106, n_542, n_370);
  nand g429 (n_543, n_368, n_369);
  nand g430 (n_544, n_370, n_369);
  nand g431 (n_545, n_368, n_370);
  nand g432 (n_88, n_543, n_544, n_545);
  xor g433 (n_371, in_2[5], in_3[5]);
  and g434 (n_380, in_2[5], in_3[5]);
  xor g435 (n_546, n_371, n_372);
  xor g436 (n_378, n_546, n_373);
  nand g437 (n_547, n_371, n_372);
  nand g438 (n_548, n_373, n_372);
  nand g439 (n_549, n_371, n_373);
  nand g440 (n_387, n_547, n_548, n_549);
  xor g441 (n_550, n_374, n_375);
  xor g442 (n_379, n_550, n_376);
  nand g443 (n_551, n_374, n_375);
  nand g444 (n_552, n_376, n_375);
  nand g445 (n_553, n_374, n_376);
  nand g446 (n_386, n_551, n_552, n_553);
  xor g447 (n_554, n_377, n_378);
  xor g448 (n_105, n_554, n_379);
  nand g449 (n_555, n_377, n_378);
  nand g450 (n_556, n_379, n_378);
  nand g451 (n_557, n_377, n_379);
  nand g452 (n_87, n_555, n_556, n_557);
  xor g453 (n_558, in_2[6], in_3[6]);
  xor g454 (n_384, n_558, n_380);
  nand g455 (n_559, in_2[6], in_3[6]);
  nand g456 (n_560, n_380, in_3[6]);
  nand g457 (n_561, in_2[6], n_380);
  nand g458 (n_392, n_559, n_560, n_561);
  xor g459 (n_562, n_381, n_382);
  xor g460 (n_388, n_562, n_383);
  nand g461 (n_563, n_381, n_382);
  nand g462 (n_564, n_383, n_382);
  nand g463 (n_565, n_381, n_383);
  nand g464 (n_398, n_563, n_564, n_565);
  xor g465 (n_566, n_384, n_385);
  xor g466 (n_389, n_566, n_386);
  nand g467 (n_567, n_384, n_385);
  nand g468 (n_568, n_386, n_385);
  nand g469 (n_569, n_384, n_386);
  nand g470 (n_400, n_567, n_568, n_569);
  xor g471 (n_570, n_387, n_388);
  xor g472 (n_104, n_570, n_389);
  nand g473 (n_571, n_387, n_388);
  nand g474 (n_572, n_389, n_388);
  nand g475 (n_573, n_387, n_389);
  nand g476 (n_86, n_571, n_572, n_573);
  xor g477 (n_390, in_2[7], in_3[7]);
  and g478 (n_402, in_2[7], in_3[7]);
  xor g479 (n_574, n_390, n_391);
  xor g480 (n_397, n_574, n_392);
  nand g481 (n_575, n_390, n_391);
  nand g482 (n_576, n_392, n_391);
  nand g483 (n_577, n_390, n_392);
  nand g484 (n_410, n_575, n_576, n_577);
  xor g485 (n_578, n_393, n_394);
  xor g486 (n_399, n_578, n_395);
  nand g487 (n_579, n_393, n_394);
  nand g488 (n_580, n_395, n_394);
  nand g489 (n_581, n_393, n_395);
  nand g490 (n_409, n_579, n_580, n_581);
  xor g491 (n_582, n_396, n_397);
  xor g492 (n_401, n_582, n_398);
  nand g493 (n_583, n_396, n_397);
  nand g494 (n_584, n_398, n_397);
  nand g495 (n_585, n_396, n_398);
  nand g496 (n_413, n_583, n_584, n_585);
  xor g497 (n_586, n_399, n_400);
  xor g498 (n_103, n_586, n_401);
  nand g499 (n_587, n_399, n_400);
  nand g500 (n_588, n_401, n_400);
  nand g501 (n_589, n_399, n_401);
  nand g502 (n_85, n_587, n_588, n_589);
  xor g503 (n_590, in_2[8], in_3[8]);
  xor g504 (n_404, n_590, n_402);
  nand g505 (n_591, in_2[8], in_3[8]);
  nand g506 (n_592, n_402, in_3[8]);
  nand g507 (n_593, in_2[8], n_402);
  nand g508 (n_417, n_591, n_592, n_593);
  xor g509 (n_594, n_403, n_404);
  xor g510 (n_411, n_594, n_405);
  nand g511 (n_595, n_403, n_404);
  nand g512 (n_596, n_405, n_404);
  nand g513 (n_597, n_403, n_405);
  nand g514 (n_423, n_595, n_596, n_597);
  xor g515 (n_598, n_406, n_407);
  xor g516 (n_412, n_598, n_408);
  nand g517 (n_599, n_406, n_407);
  nand g518 (n_600, n_408, n_407);
  nand g519 (n_601, n_406, n_408);
  nand g520 (n_422, n_599, n_600, n_601);
  xor g521 (n_602, n_409, n_410);
  xor g522 (n_414, n_602, n_411);
  nand g523 (n_603, n_409, n_410);
  nand g524 (n_604, n_411, n_410);
  nand g525 (n_605, n_409, n_411);
  nand g526 (n_427, n_603, n_604, n_605);
  xor g527 (n_606, n_412, n_413);
  xor g528 (n_102, n_606, n_414);
  nand g529 (n_607, n_412, n_413);
  nand g530 (n_608, n_414, n_413);
  nand g531 (n_609, n_412, n_414);
  nand g532 (n_84, n_607, n_608, n_609);
  xor g533 (n_610, in_2[9], in_3[9]);
  nand g535 (n_611, in_2[9], in_3[9]);
  nand g538 (n_433, n_611, n_873, n_874);
  xor g539 (n_614, n_416, n_417);
  xor g540 (n_424, n_614, n_418);
  nand g541 (n_615, n_416, n_417);
  nand g542 (n_616, n_418, n_417);
  nand g543 (n_617, n_416, n_418);
  nand g544 (n_434, n_615, n_616, n_617);
  xor g545 (n_618, n_419, n_420);
  xor g546 (n_425, n_618, n_421);
  nand g547 (n_619, n_419, n_420);
  nand g548 (n_620, n_421, n_420);
  nand g549 (n_621, n_419, n_421);
  nand g550 (n_437, n_619, n_620, n_621);
  xor g551 (n_622, n_422, n_423);
  xor g552 (n_426, n_622, n_424);
  nand g553 (n_623, n_422, n_423);
  nand g554 (n_624, n_424, n_423);
  nand g555 (n_625, n_422, n_424);
  nand g556 (n_439, n_623, n_624, n_625);
  xor g557 (n_626, n_425, n_426);
  xor g558 (n_101, n_626, n_427);
  nand g559 (n_627, n_425, n_426);
  nand g560 (n_628, n_427, n_426);
  nand g561 (n_629, n_425, n_427);
  nand g562 (n_83, n_627, n_628, n_629);
  xor g563 (n_630, in_2[10], in_3[10]);
  xor g564 (n_435, n_630, n_428);
  nand g565 (n_631, in_2[10], in_3[10]);
  nand g566 (n_632, n_428, in_3[10]);
  nand g567 (n_633, in_2[10], n_428);
  nand g568 (n_446, n_631, n_632, n_633);
  xor g569 (n_634, n_429, n_430);
  xor g570 (n_436, n_634, n_431);
  nand g571 (n_635, n_429, n_430);
  nand g572 (n_636, n_431, n_430);
  nand g573 (n_637, n_429, n_431);
  nand g574 (n_447, n_635, n_636, n_637);
  xor g576 (n_438, n_876, n_434);
  nand g578 (n_640, n_434, n_433);
  nand g580 (n_450, n_877, n_640, n_878);
  xor g581 (n_642, n_435, n_436);
  xor g582 (n_440, n_642, n_437);
  nand g583 (n_643, n_435, n_436);
  nand g584 (n_644, n_437, n_436);
  nand g585 (n_645, n_435, n_437);
  nand g586 (n_453, n_643, n_644, n_645);
  xor g587 (n_646, n_438, n_439);
  xor g588 (n_100, n_646, n_440);
  nand g589 (n_647, n_438, n_439);
  nand g590 (n_648, n_440, n_439);
  nand g591 (n_649, n_438, n_440);
  nand g592 (n_82, n_647, n_648, n_649);
  xor g593 (n_650, in_2[11], in_3[11]);
  xor g594 (n_448, n_650, n_441);
  nand g595 (n_651, in_2[11], in_3[11]);
  nand g596 (n_652, n_441, in_3[11]);
  nand g597 (n_653, in_2[11], n_441);
  nand g598 (n_459, n_651, n_652, n_653);
  xor g599 (n_654, n_442, n_443);
  xor g600 (n_449, n_654, n_444);
  nand g601 (n_655, n_442, n_443);
  nand g602 (n_656, n_444, n_443);
  nand g603 (n_657, n_442, n_444);
  nand g604 (n_460, n_655, n_656, n_657);
  xor g606 (n_451, n_879, n_447);
  nand g608 (n_660, n_447, n_446);
  nand g610 (n_463, n_880, n_660, n_881);
  xor g611 (n_662, n_448, n_449);
  xor g612 (n_452, n_662, n_450);
  nand g613 (n_663, n_448, n_449);
  nand g614 (n_664, n_450, n_449);
  nand g615 (n_665, n_448, n_450);
  nand g616 (n_466, n_663, n_664, n_665);
  xor g617 (n_666, n_451, n_452);
  xor g618 (n_99, n_666, n_453);
  nand g619 (n_667, n_451, n_452);
  nand g620 (n_668, n_453, n_452);
  nand g621 (n_669, n_451, n_453);
  nand g622 (n_81, n_667, n_668, n_669);
  xor g623 (n_670, in_2[12], in_3[12]);
  xor g624 (n_461, n_670, n_454);
  nand g625 (n_671, in_2[12], in_3[12]);
  nand g626 (n_672, n_454, in_3[12]);
  nand g627 (n_673, in_2[12], n_454);
  nand g628 (n_472, n_671, n_672, n_673);
  xor g629 (n_674, n_455, n_456);
  xor g630 (n_462, n_674, n_457);
  nand g631 (n_675, n_455, n_456);
  nand g632 (n_676, n_457, n_456);
  nand g633 (n_677, n_455, n_457);
  nand g634 (n_473, n_675, n_676, n_677);
  xor g636 (n_464, n_882, n_460);
  nand g638 (n_680, n_460, n_459);
  nand g640 (n_476, n_883, n_680, n_884);
  xor g641 (n_682, n_461, n_462);
  xor g642 (n_465, n_682, n_463);
  nand g643 (n_683, n_461, n_462);
  nand g644 (n_684, n_463, n_462);
  nand g645 (n_685, n_461, n_463);
  nand g646 (n_479, n_683, n_684, n_685);
  xor g647 (n_686, n_464, n_465);
  xor g648 (n_98, n_686, n_466);
  nand g649 (n_687, n_464, n_465);
  nand g650 (n_688, n_466, n_465);
  nand g651 (n_689, n_464, n_466);
  nand g652 (n_80, n_687, n_688, n_689);
  xor g653 (n_690, in_2[13], in_3[13]);
  xor g654 (n_474, n_690, n_467);
  nand g655 (n_691, in_2[13], in_3[13]);
  nand g656 (n_692, n_467, in_3[13]);
  nand g657 (n_693, in_2[13], n_467);
  nand g658 (n_485, n_691, n_692, n_693);
  xor g659 (n_694, n_468, n_469);
  xor g660 (n_475, n_694, n_470);
  nand g661 (n_695, n_468, n_469);
  nand g662 (n_696, n_470, n_469);
  nand g663 (n_697, n_468, n_470);
  nand g664 (n_486, n_695, n_696, n_697);
  xor g666 (n_477, n_885, n_473);
  nand g668 (n_700, n_473, n_472);
  nand g670 (n_489, n_886, n_700, n_887);
  xor g671 (n_702, n_474, n_475);
  xor g672 (n_478, n_702, n_476);
  nand g673 (n_703, n_474, n_475);
  nand g674 (n_704, n_476, n_475);
  nand g675 (n_705, n_474, n_476);
  nand g676 (n_492, n_703, n_704, n_705);
  xor g677 (n_706, n_477, n_478);
  xor g678 (n_97, n_706, n_479);
  nand g679 (n_707, n_477, n_478);
  nand g680 (n_708, n_479, n_478);
  nand g681 (n_709, n_477, n_479);
  nand g682 (n_79, n_707, n_708, n_709);
  xor g683 (n_710, in_2[14], in_3[14]);
  xor g684 (n_487, n_710, n_480);
  nand g685 (n_711, in_2[14], in_3[14]);
  nand g686 (n_712, n_480, in_3[14]);
  nand g687 (n_713, in_2[14], n_480);
  nand g688 (n_498, n_711, n_712, n_713);
  xor g689 (n_714, n_481, n_482);
  xor g690 (n_488, n_714, n_483);
  nand g691 (n_715, n_481, n_482);
  nand g692 (n_716, n_483, n_482);
  nand g693 (n_717, n_481, n_483);
  nand g694 (n_499, n_715, n_716, n_717);
  xor g696 (n_490, n_888, n_486);
  nand g698 (n_720, n_486, n_485);
  nand g700 (n_502, n_889, n_720, n_890);
  xor g701 (n_722, n_487, n_488);
  xor g702 (n_491, n_722, n_489);
  nand g703 (n_723, n_487, n_488);
  nand g704 (n_724, n_489, n_488);
  nand g705 (n_725, n_487, n_489);
  nand g706 (n_505, n_723, n_724, n_725);
  xor g707 (n_726, n_490, n_491);
  xor g708 (n_96, n_726, n_492);
  nand g709 (n_727, n_490, n_491);
  nand g710 (n_728, n_492, n_491);
  nand g711 (n_729, n_490, n_492);
  nand g712 (n_78, n_727, n_728, n_729);
  xor g713 (n_730, in_2[15], in_3[15]);
  xor g714 (n_500, n_730, n_493);
  nand g715 (n_731, in_2[15], in_3[15]);
  nand g716 (n_732, n_493, in_3[15]);
  nand g717 (n_733, in_2[15], n_493);
  nand g718 (n_512, n_731, n_732, n_733);
  xor g719 (n_734, n_494, n_495);
  xor g720 (n_501, n_734, n_496);
  nand g721 (n_735, n_494, n_495);
  nand g722 (n_736, n_496, n_495);
  nand g723 (n_737, n_494, n_496);
  nand g724 (n_511, n_735, n_736, n_737);
  xor g726 (n_503, n_891, n_499);
  nand g728 (n_740, n_499, n_498);
  nand g730 (n_514, n_892, n_740, n_893);
  xor g731 (n_742, n_500, n_501);
  xor g732 (n_504, n_742, n_502);
  nand g733 (n_743, n_500, n_501);
  nand g734 (n_744, n_502, n_501);
  nand g735 (n_745, n_500, n_502);
  nand g736 (n_517, n_743, n_744, n_745);
  xor g737 (n_746, n_503, n_504);
  xor g738 (n_95, n_746, n_505);
  nand g739 (n_747, n_503, n_504);
  nand g740 (n_748, n_505, n_504);
  nand g741 (n_749, n_503, n_505);
  nand g742 (n_77, n_747, n_748, n_749);
  xor g743 (n_750, n_506, n_507);
  xor g744 (n_513, n_750, n_508);
  xor g750 (n_515, n_875, n_511);
  xor g755 (n_758, n_512, n_513);
  xor g756 (n_516, n_758, n_514);
  xor g761 (n_762, n_515, n_516);
  xor g762 (n_94, n_762, n_517);
  xor g767 (n_864, in_3[0], n_110);
  nand g768 (n_766, in_3[0], n_110);
  nand g769 (n_767, in_3[0], in_2[0]);
  nand g770 (n_768, n_110, in_2[0]);
  nand g771 (n_770, n_766, n_767, n_768);
  nor g772 (n_769, n_92, n_109);
  nand g773 (n_772, n_92, n_109);
  nor g774 (n_774, n_91, n_108);
  nand g775 (n_777, n_91, n_108);
  nor g776 (n_779, n_90, n_107);
  nand g777 (n_782, n_90, n_107);
  nor g778 (n_784, n_89, n_106);
  nand g779 (n_787, n_89, n_106);
  nor g780 (n_789, n_88, n_105);
  nand g781 (n_792, n_88, n_105);
  nor g782 (n_794, n_87, n_104);
  nand g783 (n_797, n_87, n_104);
  nor g784 (n_799, n_86, n_103);
  nand g785 (n_802, n_86, n_103);
  nor g786 (n_804, n_85, n_102);
  nand g787 (n_807, n_85, n_102);
  nor g788 (n_809, n_84, n_101);
  nand g789 (n_812, n_84, n_101);
  nor g790 (n_814, n_83, n_100);
  nand g791 (n_817, n_83, n_100);
  nor g792 (n_819, n_82, n_99);
  nand g793 (n_822, n_82, n_99);
  nor g794 (n_824, n_81, n_98);
  nand g795 (n_827, n_81, n_98);
  nor g796 (n_829, n_80, n_97);
  nand g797 (n_832, n_80, n_97);
  nor g798 (n_834, n_79, n_96);
  nand g799 (n_837, n_79, n_96);
  nor g800 (n_839, n_78, n_95);
  nand g801 (n_842, n_78, n_95);
  nor g802 (n_844, n_77, n_94);
  nand g803 (n_847, n_77, n_94);
  nand g806 (n_775, n_772, n_894);
  nand g809 (n_780, n_777, n_897);
  nand g812 (n_785, n_782, n_900);
  nand g815 (n_790, n_787, n_903);
  nand g818 (n_795, n_792, n_910);
  nand g821 (n_800, n_797, n_915);
  nand g824 (n_805, n_802, n_916);
  nand g827 (n_810, n_807, n_917);
  nand g830 (n_815, n_812, n_918);
  nand g833 (n_820, n_817, n_919);
  nand g836 (n_825, n_822, n_920);
  nand g839 (n_830, n_827, n_921);
  nand g842 (n_835, n_832, n_922);
  nand g845 (n_840, n_837, n_923);
  nand g848 (n_845, n_842, n_924);
  xnor g851 (out_0[1], n_770, n_895);
  xnor g853 (out_0[2], n_775, n_896);
  xnor g855 (out_0[3], n_780, n_898);
  xnor g857 (out_0[4], n_785, n_899);
  xnor g859 (out_0[5], n_790, n_901);
  xnor g861 (out_0[6], n_795, n_902);
  xnor g863 (out_0[7], n_800, n_904);
  xnor g865 (out_0[8], n_805, n_905);
  xnor g867 (out_0[9], n_810, n_906);
  xnor g869 (out_0[10], n_815, n_907);
  xnor g871 (out_0[11], n_820, n_908);
  xnor g873 (out_0[12], n_825, n_909);
  xnor g875 (out_0[13], n_830, n_911);
  xnor g877 (out_0[14], n_835, n_912);
  xnor g879 (out_0[15], n_840, n_913);
  xnor g881 (out_0[16], n_845, n_914);
  xor g882 (out_0[0], in_2[0], n_864);
  and g884 (n_867, wc, n_221);
  not gc (wc, in_0[0]);
  and g885 (n_868, wc0, n_270);
  not gc0 (wc0, in_0[0]);
  and g886 (n_869, wc1, n_313);
  not gc1 (wc1, in_0[0]);
  and g887 (n_117, wc2, n_115);
  not gc2 (wc2, in_1[0]);
  and g889 (n_176, n_174, wc3);
  not gc3 (wc3, n_172);
  and g890 (n_229, n_227, wc4);
  not gc4 (wc4, n_225);
  and g891 (n_278, n_276, wc5);
  not gc5 (wc5, n_274);
  and g892 (n_354, in_1[1], wc6);
  not gc6 (wc6, n_110);
  xnor g901 (n_421, n_326, n_610);
  or g902 (n_873, wc7, n_326);
  not gc7 (wc7, in_3[9]);
  or g903 (n_874, wc8, n_326);
  not gc8 (wc8, in_2[9]);
  xnor g904 (n_875, n_510, n_347);
  xnor g905 (n_876, n_329, n_433);
  or g906 (n_877, wc9, n_329);
  not gc9 (wc9, n_433);
  or g907 (n_878, wc10, n_329);
  not gc10 (wc10, n_434);
  xnor g908 (n_879, n_332, n_446);
  or g909 (n_880, wc11, n_332);
  not gc11 (wc11, n_446);
  or g910 (n_881, wc12, n_332);
  not gc12 (wc12, n_447);
  xnor g911 (n_882, n_335, n_459);
  or g912 (n_883, wc13, n_335);
  not gc13 (wc13, n_459);
  or g913 (n_884, wc14, n_335);
  not gc14 (wc14, n_460);
  xnor g914 (n_885, n_338, n_472);
  or g915 (n_886, wc15, n_338);
  not gc15 (wc15, n_472);
  or g916 (n_887, wc16, n_338);
  not gc16 (wc16, n_473);
  xnor g917 (n_888, n_341, n_485);
  or g918 (n_889, wc17, n_341);
  not gc17 (wc17, n_485);
  or g919 (n_890, wc18, n_341);
  not gc18 (wc18, n_486);
  xnor g920 (n_891, n_344, n_498);
  or g921 (n_892, wc19, n_344);
  not gc19 (wc19, n_498);
  or g922 (n_893, wc20, n_344);
  not gc20 (wc20, n_499);
  or g923 (n_894, n_769, wc21);
  not gc21 (wc21, n_770);
  or g924 (n_895, wc22, n_769);
  not gc22 (wc22, n_772);
  or g925 (n_896, wc23, n_774);
  not gc23 (wc23, n_777);
  or g926 (n_897, wc24, n_774);
  not gc24 (wc24, n_775);
  or g927 (n_898, wc25, n_779);
  not gc25 (wc25, n_782);
  or g928 (n_899, wc26, n_784);
  not gc26 (wc26, n_787);
  or g929 (n_900, wc27, n_779);
  not gc27 (wc27, n_780);
  or g930 (n_901, wc28, n_789);
  not gc28 (wc28, n_792);
  or g931 (n_902, wc29, n_794);
  not gc29 (wc29, n_797);
  or g932 (n_903, wc30, n_784);
  not gc30 (wc30, n_785);
  or g933 (n_904, wc31, n_799);
  not gc31 (wc31, n_802);
  or g934 (n_905, wc32, n_804);
  not gc32 (wc32, n_807);
  or g935 (n_906, wc33, n_809);
  not gc33 (wc33, n_812);
  or g936 (n_907, wc34, n_814);
  not gc34 (wc34, n_817);
  or g937 (n_908, wc35, n_819);
  not gc35 (wc35, n_822);
  or g938 (n_909, wc36, n_824);
  not gc36 (wc36, n_827);
  or g939 (n_910, wc37, n_789);
  not gc37 (wc37, n_790);
  or g940 (n_911, wc38, n_829);
  not gc38 (wc38, n_832);
  or g941 (n_912, wc39, n_834);
  not gc39 (wc39, n_837);
  or g942 (n_913, wc40, n_839);
  not gc40 (wc40, n_842);
  or g943 (n_914, wc41, n_844);
  not gc41 (wc41, n_847);
  or g944 (n_915, wc42, n_794);
  not gc42 (wc42, n_795);
  or g945 (n_916, wc43, n_799);
  not gc43 (wc43, n_800);
  or g946 (n_917, wc44, n_804);
  not gc44 (wc44, n_805);
  or g947 (n_918, wc45, n_809);
  not gc45 (wc45, n_810);
  or g948 (n_919, wc46, n_814);
  not gc46 (wc46, n_815);
  or g949 (n_920, wc47, n_819);
  not gc47 (wc47, n_820);
  or g950 (n_921, wc48, n_824);
  not gc48 (wc48, n_825);
  or g951 (n_922, wc49, n_829);
  not gc49 (wc49, n_830);
  or g952 (n_923, wc50, n_834);
  not gc50 (wc50, n_835);
  or g953 (n_924, wc51, n_839);
  not gc51 (wc51, n_840);
endmodule

module csa_tree_add_25_30_group_50_GENERIC(in_0, in_1, in_2, in_3,
     out_0);
  input [16:0] in_0, in_2, in_3;
  input [7:0] in_1;
  output [16:0] out_0;
  wire [16:0] in_0, in_2, in_3;
  wire [7:0] in_1;
  wire [16:0] out_0;
  csa_tree_add_25_30_group_50_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .out_0 (out_0));
endmodule

module csa_tree_mul_25_40_group_52_GENERIC_REAL(in_0, in_1, out_0);
// synthesis_equation "assign out_0 = ( in_0 * in_1 )  ;"
  input [15:0] in_0;
  input [7:0] in_1;
  output [16:0] out_0;
  wire [15:0] in_0;
  wire [7:0] in_1;
  wire [16:0] out_0;
  wire n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_79, n_80, n_81, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_131, n_137, n_139, n_140, n_141, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_188, n_190, n_191, n_192, n_194, n_195, n_196, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_237, n_239, n_240, n_241, n_243;
  wire n_244, n_245, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_280, n_282, n_283, n_293, n_296, n_299, n_302, n_305;
  wire n_308, n_311, n_314, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_355, n_356, n_358, n_359;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_369;
  wire n_370, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_387, n_388;
  wire n_389, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_399, n_400, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_493, n_497, n_498;
  wire n_499, n_500, n_501, n_505, n_506, n_507, n_508, n_509;
  wire n_510, n_511, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_529, n_530, n_531, n_532, n_533;
  wire n_534, n_535, n_536, n_537, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_553, n_554, n_555;
  wire n_556, n_557, n_558, n_559, n_560, n_561, n_566, n_570;
  wire n_577, n_580, n_582, n_585, n_587, n_588, n_590, n_592;
  wire n_593, n_595, n_597, n_598, n_600, n_602, n_603, n_605;
  wire n_607, n_608, n_610, n_612, n_613, n_615, n_617, n_618;
  wire n_620, n_622, n_623, n_625, n_627, n_628, n_630, n_632;
  wire n_633, n_635, n_637, n_638, n_640, n_642, n_643, n_645;
  wire n_647, n_648, n_650, n_652, n_653, n_655, n_676, n_677;
  wire n_678, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696;
  wire n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_705;
  wire n_706, n_708, n_709, n_710, n_711, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738;
  xor g2 (n_79, in_1[1], in_1[0]);
  xor g8 (n_80, in_1[1], in_0[0]);
  and g12 (out_0[0], in_0[0], in_1[0]);
  xor g13 (n_85, in_1[1], in_0[1]);
  nand g14 (n_86, n_85, in_1[0]);
  nand g15 (n_87, n_80, n_81);
  nand g16 (n_74, n_86, n_87);
  xor g17 (n_88, in_1[1], in_0[2]);
  nand g18 (n_89, n_88, in_1[0]);
  nand g19 (n_90, n_85, n_81);
  nand g20 (n_73, n_89, n_90);
  xor g21 (n_91, in_1[1], in_0[3]);
  nand g22 (n_92, n_91, in_1[0]);
  nand g23 (n_93, n_88, n_81);
  nand g24 (n_322, n_92, n_93);
  xor g25 (n_94, in_1[1], in_0[4]);
  nand g26 (n_95, n_94, in_1[0]);
  nand g27 (n_96, n_91, n_81);
  nand g28 (n_325, n_95, n_96);
  xor g29 (n_97, in_1[1], in_0[5]);
  nand g30 (n_98, n_97, in_1[0]);
  nand g31 (n_99, n_94, n_81);
  nand g32 (n_327, n_98, n_99);
  xor g33 (n_100, in_1[1], in_0[6]);
  nand g34 (n_101, n_100, in_1[0]);
  nand g35 (n_102, n_97, n_81);
  nand g36 (n_332, n_101, n_102);
  xor g37 (n_103, in_1[1], in_0[7]);
  nand g38 (n_104, n_103, in_1[0]);
  nand g39 (n_105, n_100, n_81);
  nand g40 (n_338, n_104, n_105);
  xor g41 (n_106, in_1[1], in_0[8]);
  nand g42 (n_107, n_106, in_1[0]);
  nand g43 (n_108, n_103, n_81);
  nand g44 (n_346, n_107, n_108);
  xor g45 (n_109, in_1[1], in_0[9]);
  nand g46 (n_110, n_109, in_1[0]);
  nand g47 (n_111, n_106, n_81);
  nand g48 (n_358, n_110, n_111);
  xor g49 (n_112, in_1[1], in_0[10]);
  nand g50 (n_113, n_112, in_1[0]);
  nand g51 (n_114, n_109, n_81);
  nand g52 (n_365, n_113, n_114);
  xor g53 (n_115, in_1[1], in_0[11]);
  nand g54 (n_116, n_115, in_1[0]);
  nand g55 (n_117, n_112, n_81);
  nand g56 (n_376, n_116, n_117);
  xor g57 (n_118, in_1[1], in_0[12]);
  nand g58 (n_119, n_118, in_1[0]);
  nand g59 (n_120, n_115, n_81);
  nand g60 (n_387, n_119, n_120);
  xor g61 (n_121, in_1[1], in_0[13]);
  nand g62 (n_122, n_121, in_1[0]);
  nand g63 (n_123, n_118, n_81);
  nand g64 (n_398, n_122, n_123);
  xor g65 (n_124, in_1[1], in_0[14]);
  nand g66 (n_125, n_124, in_1[0]);
  nand g67 (n_126, n_121, n_81);
  nand g68 (n_409, n_125, n_126);
  xor g69 (n_127, in_1[1], in_0[15]);
  nand g70 (n_128, n_127, in_1[0]);
  nand g71 (n_129, n_124, n_81);
  nand g72 (n_420, n_128, n_129);
  nand g74 (n_131, in_1[1], in_1[0]);
  nand g75 (n_75, n_127, n_81);
  nand g76 (n_431, n_131, n_75);
  xor g81 (n_137, in_1[2], in_1[1]);
  xor g82 (n_139, in_1[3], in_1[2]);
  nor g86 (n_190, in_1[1], in_1[2]);
  nand g87 (n_188, in_1[1], in_1[2]);
  xor g88 (n_140, in_1[3], in_0[0]);
  and g92 (n_56, in_0[0], n_137);
  xor g93 (n_145, in_1[3], in_0[1]);
  nand g94 (n_146, n_145, n_137);
  nand g95 (n_147, n_140, n_141);
  nand g96 (n_55, n_146, n_147);
  xor g97 (n_148, in_1[3], in_0[2]);
  nand g98 (n_149, n_148, n_137);
  nand g99 (n_150, n_145, n_141);
  nand g100 (n_324, n_149, n_150);
  xor g101 (n_151, in_1[3], in_0[3]);
  nand g102 (n_152, n_151, n_137);
  nand g103 (n_153, n_148, n_141);
  nand g104 (n_328, n_152, n_153);
  xor g105 (n_154, in_1[3], in_0[4]);
  nand g106 (n_155, n_154, n_137);
  nand g107 (n_156, n_151, n_141);
  nand g108 (n_333, n_155, n_156);
  xor g109 (n_157, in_1[3], in_0[5]);
  nand g110 (n_158, n_157, n_137);
  nand g111 (n_159, n_154, n_141);
  nand g112 (n_340, n_158, n_159);
  xor g113 (n_160, in_1[3], in_0[6]);
  nand g114 (n_161, n_160, n_137);
  nand g115 (n_162, n_157, n_141);
  nand g116 (n_348, n_161, n_162);
  xor g117 (n_163, in_1[3], in_0[7]);
  nand g118 (n_164, n_163, n_137);
  nand g119 (n_165, n_160, n_141);
  nand g120 (n_355, n_164, n_165);
  xor g121 (n_166, in_1[3], in_0[8]);
  nand g122 (n_167, n_166, n_137);
  nand g123 (n_168, n_163, n_141);
  nand g124 (n_366, n_167, n_168);
  xor g125 (n_169, in_1[3], in_0[9]);
  nand g126 (n_170, n_169, n_137);
  nand g127 (n_171, n_166, n_141);
  nand g128 (n_377, n_170, n_171);
  xor g129 (n_172, in_1[3], in_0[10]);
  nand g130 (n_173, n_172, n_137);
  nand g131 (n_174, n_169, n_141);
  nand g132 (n_388, n_173, n_174);
  xor g133 (n_175, in_1[3], in_0[11]);
  nand g134 (n_176, n_175, n_137);
  nand g135 (n_177, n_172, n_141);
  nand g136 (n_399, n_176, n_177);
  xor g137 (n_178, in_1[3], in_0[12]);
  nand g138 (n_179, n_178, n_137);
  nand g139 (n_180, n_175, n_141);
  nand g140 (n_410, n_179, n_180);
  xor g141 (n_181, in_1[3], in_0[13]);
  nand g142 (n_182, n_181, n_137);
  nand g143 (n_183, n_178, n_141);
  nand g144 (n_421, n_182, n_183);
  xor g145 (n_184, in_1[3], in_0[14]);
  nand g146 (n_185, n_184, n_137);
  nand g147 (n_186, n_181, n_141);
  nand g148 (n_432, n_185, n_186);
  or g151 (n_191, n_676, n_190);
  and g152 (n_321, in_1[3], n_191);
  xor g153 (n_192, in_1[4], in_1[3]);
  xor g154 (n_194, in_1[5], in_1[4]);
  nor g158 (n_239, in_1[3], in_1[4]);
  nand g159 (n_237, in_1[3], in_1[4]);
  xor g160 (n_195, in_1[5], in_0[0]);
  and g164 (n_323, in_0[0], n_192);
  xor g165 (n_200, in_1[5], in_0[1]);
  nand g166 (n_201, n_200, n_192);
  nand g167 (n_202, n_195, n_196);
  nand g168 (n_329, n_201, n_202);
  xor g169 (n_203, in_1[5], in_0[2]);
  nand g170 (n_204, n_203, n_192);
  nand g171 (n_205, n_200, n_196);
  nand g172 (n_334, n_204, n_205);
  xor g173 (n_206, in_1[5], in_0[3]);
  nand g174 (n_207, n_206, n_192);
  nand g175 (n_208, n_203, n_196);
  nand g176 (n_341, n_207, n_208);
  xor g177 (n_209, in_1[5], in_0[4]);
  nand g178 (n_210, n_209, n_192);
  nand g179 (n_211, n_206, n_196);
  nand g180 (n_349, n_210, n_211);
  xor g181 (n_212, in_1[5], in_0[5]);
  nand g182 (n_213, n_212, n_192);
  nand g183 (n_214, n_209, n_196);
  nand g184 (n_359, n_213, n_214);
  xor g185 (n_215, in_1[5], in_0[6]);
  nand g186 (n_216, n_215, n_192);
  nand g187 (n_217, n_212, n_196);
  nand g188 (n_369, n_216, n_217);
  xor g189 (n_218, in_1[5], in_0[7]);
  nand g190 (n_219, n_218, n_192);
  nand g191 (n_220, n_215, n_196);
  nand g192 (n_380, n_219, n_220);
  xor g193 (n_221, in_1[5], in_0[8]);
  nand g194 (n_222, n_221, n_192);
  nand g195 (n_223, n_218, n_196);
  nand g196 (n_391, n_222, n_223);
  xor g197 (n_224, in_1[5], in_0[9]);
  nand g198 (n_225, n_224, n_192);
  nand g199 (n_226, n_221, n_196);
  nand g200 (n_402, n_225, n_226);
  xor g201 (n_227, in_1[5], in_0[10]);
  nand g202 (n_228, n_227, n_192);
  nand g203 (n_229, n_224, n_196);
  nand g204 (n_413, n_228, n_229);
  xor g205 (n_230, in_1[5], in_0[11]);
  nand g206 (n_231, n_230, n_192);
  nand g207 (n_232, n_227, n_196);
  nand g208 (n_424, n_231, n_232);
  xor g209 (n_233, in_1[5], in_0[12]);
  nand g210 (n_234, n_233, n_192);
  nand g211 (n_235, n_230, n_196);
  nand g212 (n_435, n_234, n_235);
  or g215 (n_240, n_677, n_239);
  and g216 (n_326, in_1[5], n_240);
  xor g217 (n_241, in_1[6], in_1[5]);
  xor g218 (n_243, in_1[7], in_1[6]);
  nor g222 (n_282, in_1[5], in_1[6]);
  nand g223 (n_280, in_1[5], in_1[6]);
  xor g224 (n_244, in_1[7], in_0[0]);
  and g228 (n_331, in_0[0], n_241);
  xor g229 (n_249, in_1[7], in_0[1]);
  nand g230 (n_250, n_249, n_241);
  nand g231 (n_251, n_244, n_245);
  nand g232 (n_339, n_250, n_251);
  xor g233 (n_252, in_1[7], in_0[2]);
  nand g234 (n_253, n_252, n_241);
  nand g235 (n_254, n_249, n_245);
  nand g236 (n_347, n_253, n_254);
  xor g237 (n_255, in_1[7], in_0[3]);
  nand g238 (n_256, n_255, n_241);
  nand g239 (n_257, n_252, n_245);
  nand g240 (n_356, n_256, n_257);
  xor g241 (n_258, in_1[7], in_0[4]);
  nand g242 (n_259, n_258, n_241);
  nand g243 (n_260, n_255, n_245);
  nand g244 (n_367, n_259, n_260);
  xor g245 (n_261, in_1[7], in_0[5]);
  nand g246 (n_262, n_261, n_241);
  nand g247 (n_263, n_258, n_245);
  nand g248 (n_378, n_262, n_263);
  xor g249 (n_264, in_1[7], in_0[6]);
  nand g250 (n_265, n_264, n_241);
  nand g251 (n_266, n_261, n_245);
  nand g252 (n_389, n_265, n_266);
  xor g253 (n_267, in_1[7], in_0[7]);
  nand g254 (n_268, n_267, n_241);
  nand g255 (n_269, n_264, n_245);
  nand g256 (n_400, n_268, n_269);
  xor g257 (n_270, in_1[7], in_0[8]);
  nand g258 (n_271, n_270, n_241);
  nand g259 (n_272, n_267, n_245);
  nand g260 (n_411, n_271, n_272);
  xor g261 (n_273, in_1[7], in_0[9]);
  nand g262 (n_274, n_273, n_241);
  nand g263 (n_275, n_270, n_245);
  nand g264 (n_422, n_274, n_275);
  xor g265 (n_276, in_1[7], in_0[10]);
  nand g266 (n_277, n_276, n_241);
  nand g267 (n_278, n_273, n_245);
  nand g268 (n_433, n_277, n_278);
  or g271 (n_283, n_678, n_282);
  and g272 (n_337, in_1[7], n_283);
  and g284 (n_345, in_0[0], in_1[7]);
  nand g286 (n_293, in_0[1], in_1[7]);
  nand g290 (n_296, in_0[2], in_1[7]);
  nand g294 (n_299, in_0[3], in_1[7]);
  nand g298 (n_302, in_0[4], in_1[7]);
  nand g302 (n_305, in_0[5], in_1[7]);
  nand g306 (n_308, in_0[6], in_1[7]);
  nand g310 (n_311, in_0[7], in_1[7]);
  nand g314 (n_314, in_0[8], in_1[7]);
  xor g365 (n_72, n_321, n_322);
  and g366 (n_54, n_321, n_322);
  xor g367 (n_442, n_323, n_324);
  xor g368 (n_71, n_442, n_325);
  nand g369 (n_443, n_323, n_324);
  nand g370 (n_444, n_325, n_324);
  nand g371 (n_445, n_323, n_325);
  nand g372 (n_53, n_443, n_444, n_445);
  xor g373 (n_330, n_326, n_327);
  and g374 (n_335, n_326, n_327);
  xor g375 (n_446, n_328, n_329);
  xor g376 (n_70, n_446, n_330);
  nand g377 (n_447, n_328, n_329);
  nand g378 (n_448, n_330, n_329);
  nand g379 (n_449, n_328, n_330);
  nand g380 (n_52, n_447, n_448, n_449);
  xor g381 (n_450, n_331, n_332);
  xor g382 (n_336, n_450, n_333);
  nand g383 (n_451, n_331, n_332);
  nand g384 (n_452, n_333, n_332);
  nand g385 (n_453, n_331, n_333);
  nand g386 (n_343, n_451, n_452, n_453);
  xor g387 (n_454, n_334, n_335);
  xor g388 (n_69, n_454, n_336);
  nand g389 (n_455, n_334, n_335);
  nand g390 (n_456, n_336, n_335);
  nand g391 (n_457, n_334, n_336);
  nand g392 (n_51, n_455, n_456, n_457);
  xor g393 (n_342, n_337, n_338);
  and g394 (n_350, n_337, n_338);
  xor g395 (n_458, n_339, n_340);
  xor g396 (n_344, n_458, n_341);
  nand g397 (n_459, n_339, n_340);
  nand g398 (n_460, n_341, n_340);
  nand g399 (n_461, n_339, n_341);
  nand g400 (n_351, n_459, n_460, n_461);
  xor g401 (n_462, n_342, n_343);
  xor g402 (n_68, n_462, n_344);
  nand g403 (n_463, n_342, n_343);
  nand g404 (n_464, n_344, n_343);
  nand g405 (n_465, n_342, n_344);
  nand g406 (n_50, n_463, n_464, n_465);
  xor g407 (n_466, n_345, n_346);
  xor g408 (n_352, n_466, n_347);
  nand g409 (n_467, n_345, n_346);
  nand g410 (n_468, n_347, n_346);
  nand g411 (n_469, n_345, n_347);
  nand g412 (n_361, n_467, n_468, n_469);
  xor g413 (n_470, n_348, n_349);
  xor g414 (n_353, n_470, n_350);
  nand g415 (n_471, n_348, n_349);
  nand g416 (n_472, n_350, n_349);
  nand g417 (n_473, n_348, n_350);
  nand g418 (n_363, n_471, n_472, n_473);
  xor g419 (n_474, n_351, n_352);
  xor g420 (n_67, n_474, n_353);
  nand g421 (n_475, n_351, n_352);
  nand g422 (n_476, n_353, n_352);
  nand g423 (n_477, n_351, n_353);
  nand g424 (n_49, n_475, n_476, n_477);
  xor g428 (n_362, n_682, n_358);
  nand g431 (n_481, n_356, n_358);
  nand g432 (n_372, n_683, n_684, n_481);
  xor g433 (n_482, n_359, n_355);
  xor g434 (n_364, n_482, n_361);
  nand g435 (n_483, n_359, n_355);
  nand g436 (n_484, n_361, n_355);
  nand g437 (n_485, n_359, n_361);
  nand g438 (n_375, n_483, n_484, n_485);
  xor g439 (n_486, n_362, n_363);
  xor g440 (n_66, n_486, n_364);
  nand g441 (n_487, n_362, n_363);
  nand g442 (n_488, n_364, n_363);
  nand g443 (n_489, n_362, n_364);
  nand g444 (n_48, n_487, n_488, n_489);
  xor g445 (n_370, n_365, n_366);
  and g446 (n_382, n_365, n_366);
  xor g448 (n_373, n_685, n_369);
  nand g451 (n_493, n_367, n_369);
  nand g452 (n_383, n_686, n_687, n_493);
  xor g454 (n_374, n_370, n_372);
  nand g457 (n_497, n_370, n_372);
  xor g459 (n_498, n_373, n_374);
  xor g460 (n_65, n_498, n_375);
  nand g461 (n_499, n_373, n_374);
  nand g462 (n_500, n_375, n_374);
  nand g463 (n_501, n_373, n_375);
  nand g464 (n_47, n_499, n_500, n_501);
  xor g465 (n_381, n_376, n_377);
  and g466 (n_393, n_376, n_377);
  xor g468 (n_384, n_688, n_380);
  nand g471 (n_505, n_378, n_380);
  nand g472 (n_394, n_689, n_690, n_505);
  xor g473 (n_506, n_381, n_382);
  xor g474 (n_385, n_506, n_383);
  nand g475 (n_507, n_381, n_382);
  nand g476 (n_508, n_383, n_382);
  nand g477 (n_509, n_381, n_383);
  nand g478 (n_397, n_507, n_508, n_509);
  xor g479 (n_510, n_384, n_385);
  nand g481 (n_511, n_384, n_385);
  nand g484 (n_46, n_511, n_709, n_710);
  xor g485 (n_392, n_387, n_388);
  and g486 (n_404, n_387, n_388);
  xor g488 (n_395, n_691, n_391);
  nand g491 (n_517, n_389, n_391);
  nand g492 (n_405, n_692, n_693, n_517);
  xor g493 (n_518, n_392, n_393);
  xor g494 (n_396, n_518, n_394);
  nand g495 (n_519, n_392, n_393);
  nand g496 (n_520, n_394, n_393);
  nand g497 (n_521, n_392, n_394);
  nand g498 (n_408, n_519, n_520, n_521);
  xor g499 (n_522, n_395, n_396);
  xor g500 (n_63, n_522, n_397);
  nand g501 (n_523, n_395, n_396);
  nand g502 (n_524, n_397, n_396);
  nand g503 (n_525, n_395, n_397);
  nand g504 (n_45, n_523, n_524, n_525);
  xor g505 (n_403, n_398, n_399);
  and g506 (n_415, n_398, n_399);
  xor g508 (n_406, n_694, n_402);
  nand g511 (n_529, n_400, n_402);
  nand g512 (n_416, n_695, n_696, n_529);
  xor g513 (n_530, n_403, n_404);
  xor g514 (n_407, n_530, n_405);
  nand g515 (n_531, n_403, n_404);
  nand g516 (n_532, n_405, n_404);
  nand g517 (n_533, n_403, n_405);
  nand g518 (n_419, n_531, n_532, n_533);
  xor g519 (n_534, n_406, n_407);
  xor g520 (n_62, n_534, n_408);
  nand g521 (n_535, n_406, n_407);
  nand g522 (n_536, n_408, n_407);
  nand g523 (n_537, n_406, n_408);
  nand g524 (n_44, n_535, n_536, n_537);
  xor g525 (n_414, n_409, n_410);
  and g526 (n_426, n_409, n_410);
  xor g528 (n_417, n_697, n_413);
  nand g531 (n_541, n_411, n_413);
  nand g532 (n_427, n_698, n_699, n_541);
  xor g533 (n_542, n_414, n_415);
  xor g534 (n_418, n_542, n_416);
  nand g535 (n_543, n_414, n_415);
  nand g536 (n_544, n_416, n_415);
  nand g537 (n_545, n_414, n_416);
  nand g538 (n_430, n_543, n_544, n_545);
  xor g539 (n_546, n_417, n_418);
  xor g540 (n_61, n_546, n_419);
  nand g541 (n_547, n_417, n_418);
  nand g542 (n_548, n_419, n_418);
  nand g543 (n_549, n_417, n_419);
  nand g544 (n_43, n_547, n_548, n_549);
  xor g545 (n_425, n_420, n_421);
  and g546 (n_437, n_420, n_421);
  xor g548 (n_428, n_700, n_424);
  nand g551 (n_553, n_422, n_424);
  nand g552 (n_438, n_701, n_702, n_553);
  xor g553 (n_554, n_425, n_426);
  xor g554 (n_429, n_554, n_427);
  nand g555 (n_555, n_425, n_426);
  nand g556 (n_556, n_427, n_426);
  nand g557 (n_557, n_425, n_427);
  nand g558 (n_441, n_555, n_556, n_557);
  xor g559 (n_558, n_428, n_429);
  xor g560 (n_60, n_558, n_430);
  nand g561 (n_559, n_428, n_429);
  nand g562 (n_560, n_430, n_429);
  nand g563 (n_561, n_428, n_430);
  nand g564 (n_42, n_559, n_560, n_561);
  xor g565 (n_436, n_431, n_432);
  xor g568 (n_439, n_703, n_435);
  xor g573 (n_566, n_436, n_437);
  xor g574 (n_440, n_566, n_438);
  xor g579 (n_570, n_439, n_440);
  xor g580 (n_59, n_570, n_441);
  nor g590 (n_577, n_57, n_74);
  nand g591 (n_580, n_57, n_74);
  nor g592 (n_582, n_56, n_73);
  nand g593 (n_585, n_56, n_73);
  nor g594 (n_587, n_55, n_72);
  nand g595 (n_590, n_55, n_72);
  nor g596 (n_592, n_54, n_71);
  nand g597 (n_595, n_54, n_71);
  nor g598 (n_597, n_53, n_70);
  nand g599 (n_600, n_53, n_70);
  nor g600 (n_602, n_52, n_69);
  nand g601 (n_605, n_52, n_69);
  nor g602 (n_607, n_51, n_68);
  nand g603 (n_610, n_51, n_68);
  nor g604 (n_612, n_50, n_67);
  nand g605 (n_615, n_50, n_67);
  nor g606 (n_617, n_49, n_66);
  nand g607 (n_620, n_49, n_66);
  nor g608 (n_622, n_48, n_65);
  nand g609 (n_625, n_48, n_65);
  nor g610 (n_627, n_47, n_64);
  nand g611 (n_630, n_47, n_64);
  nor g612 (n_632, n_46, n_63);
  nand g613 (n_635, n_46, n_63);
  nor g614 (n_637, n_45, n_62);
  nand g615 (n_640, n_45, n_62);
  nor g616 (n_642, n_44, n_61);
  nand g617 (n_645, n_44, n_61);
  nor g618 (n_647, n_43, n_60);
  nand g619 (n_650, n_43, n_60);
  nor g620 (n_652, n_42, n_59);
  nand g621 (n_655, n_42, n_59);
  nand g627 (n_588, n_585, n_711);
  nand g630 (n_593, n_590, n_716);
  nand g633 (n_598, n_595, n_721);
  nand g636 (n_603, n_600, n_728);
  nand g639 (n_608, n_605, n_729);
  nand g642 (n_613, n_610, n_730);
  nand g645 (n_618, n_615, n_731);
  nand g648 (n_623, n_620, n_732);
  nand g651 (n_628, n_625, n_733);
  nand g654 (n_633, n_630, n_734);
  nand g657 (n_638, n_635, n_735);
  nand g660 (n_643, n_640, n_736);
  nand g663 (n_648, n_645, n_737);
  nand g666 (n_653, n_650, n_738);
  xnor g673 (out_0[3], n_588, n_708);
  xnor g675 (out_0[4], n_593, n_713);
  xnor g677 (out_0[5], n_598, n_714);
  xnor g679 (out_0[6], n_603, n_715);
  xnor g681 (out_0[7], n_608, n_717);
  xnor g683 (out_0[8], n_613, n_718);
  xnor g685 (out_0[9], n_618, n_719);
  xnor g687 (out_0[10], n_623, n_720);
  xnor g689 (out_0[11], n_628, n_722);
  xnor g691 (out_0[12], n_633, n_723);
  xnor g693 (out_0[13], n_638, n_724);
  xnor g695 (out_0[14], n_643, n_725);
  xnor g697 (out_0[15], n_648, n_726);
  xnor g699 (out_0[16], n_653, n_727);
  and g703 (n_676, wc, n_188);
  not gc (wc, in_0[0]);
  and g704 (n_677, wc0, n_237);
  not gc0 (wc0, in_0[0]);
  and g705 (n_678, wc1, n_280);
  not gc1 (wc1, in_0[0]);
  and g706 (n_81, wc2, n_79);
  not gc2 (wc2, in_1[0]);
  and g708 (n_141, n_139, wc3);
  not gc3 (wc3, n_137);
  and g709 (n_196, n_194, wc4);
  not gc4 (wc4, n_192);
  and g710 (n_245, n_243, wc5);
  not gc5 (wc5, n_241);
  and g712 (n_57, in_1[1], wc6);
  not gc6 (wc6, out_0[0]);
  xnor g721 (n_682, n_356, n_293);
  or g722 (n_683, n_293, wc7);
  not gc7 (wc7, n_356);
  or g723 (n_684, n_293, wc8);
  not gc8 (wc8, n_358);
  xnor g724 (n_685, n_367, n_296);
  or g725 (n_686, n_296, wc9);
  not gc9 (wc9, n_367);
  or g726 (n_687, n_296, wc10);
  not gc10 (wc10, n_369);
  xnor g727 (n_688, n_378, n_299);
  or g728 (n_689, n_299, wc11);
  not gc11 (wc11, n_378);
  or g729 (n_690, n_299, wc12);
  not gc12 (wc12, n_380);
  xnor g730 (n_691, n_389, n_302);
  or g731 (n_692, n_302, wc13);
  not gc13 (wc13, n_389);
  or g732 (n_693, n_302, wc14);
  not gc14 (wc14, n_391);
  xnor g733 (n_694, n_400, n_305);
  or g734 (n_695, n_305, wc15);
  not gc15 (wc15, n_400);
  or g735 (n_696, n_305, wc16);
  not gc16 (wc16, n_402);
  xnor g736 (n_697, n_411, n_308);
  or g737 (n_698, n_308, wc17);
  not gc17 (wc17, n_411);
  or g738 (n_699, n_308, wc18);
  not gc18 (wc18, n_413);
  xnor g739 (n_700, n_422, n_311);
  or g740 (n_701, n_311, wc19);
  not gc19 (wc19, n_422);
  or g741 (n_702, n_311, wc20);
  not gc20 (wc20, n_424);
  xnor g742 (n_703, n_433, n_314);
  or g743 (n_705, wc21, n_577);
  not gc21 (wc21, n_580);
  or g744 (n_706, wc22, n_582);
  not gc22 (wc22, n_585);
  not g747 (out_0[1], n_705);
  or g748 (n_708, wc23, n_587);
  not gc23 (wc23, n_590);
  xnor g749 (n_64, n_497, n_510);
  or g750 (n_709, wc24, n_497);
  not gc24 (wc24, n_385);
  or g751 (n_710, wc25, n_497);
  not gc25 (wc25, n_384);
  or g752 (n_711, n_580, n_582);
  xor g753 (out_0[2], n_580, n_706);
  or g754 (n_713, wc26, n_592);
  not gc26 (wc26, n_595);
  or g755 (n_714, wc27, n_597);
  not gc27 (wc27, n_600);
  or g756 (n_715, wc28, n_602);
  not gc28 (wc28, n_605);
  or g757 (n_716, wc29, n_587);
  not gc29 (wc29, n_588);
  or g758 (n_717, wc30, n_607);
  not gc30 (wc30, n_610);
  or g759 (n_718, wc31, n_612);
  not gc31 (wc31, n_615);
  or g760 (n_719, wc32, n_617);
  not gc32 (wc32, n_620);
  or g761 (n_720, wc33, n_622);
  not gc33 (wc33, n_625);
  or g762 (n_721, wc34, n_592);
  not gc34 (wc34, n_593);
  or g763 (n_722, wc35, n_627);
  not gc35 (wc35, n_630);
  or g764 (n_723, wc36, n_632);
  not gc36 (wc36, n_635);
  or g765 (n_724, wc37, n_637);
  not gc37 (wc37, n_640);
  or g766 (n_725, wc38, n_642);
  not gc38 (wc38, n_645);
  or g767 (n_726, wc39, n_647);
  not gc39 (wc39, n_650);
  or g768 (n_727, wc40, n_652);
  not gc40 (wc40, n_655);
  or g769 (n_728, wc41, n_597);
  not gc41 (wc41, n_598);
  or g770 (n_729, wc42, n_602);
  not gc42 (wc42, n_603);
  or g771 (n_730, wc43, n_607);
  not gc43 (wc43, n_608);
  or g772 (n_731, wc44, n_612);
  not gc44 (wc44, n_613);
  or g773 (n_732, wc45, n_617);
  not gc45 (wc45, n_618);
  or g774 (n_733, wc46, n_622);
  not gc46 (wc46, n_623);
  or g775 (n_734, wc47, n_627);
  not gc47 (wc47, n_628);
  or g776 (n_735, wc48, n_632);
  not gc48 (wc48, n_633);
  or g777 (n_736, wc49, n_637);
  not gc49 (wc49, n_638);
  or g778 (n_737, wc50, n_642);
  not gc50 (wc50, n_643);
  or g779 (n_738, wc51, n_647);
  not gc51 (wc51, n_648);
endmodule

module csa_tree_mul_25_40_group_52_GENERIC(in_0, in_1, out_0);
  input [15:0] in_0;
  input [7:0] in_1;
  output [16:0] out_0;
  wire [15:0] in_0;
  wire [7:0] in_1;
  wire [16:0] out_0;
  csa_tree_mul_25_40_group_52_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .out_0 (out_0));
endmodule

module mult_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $unsigned(A) * $unsigned(B);"
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_325;
  wire n_328, n_330, n_333, n_335, n_336, n_338, n_340, n_341;
  wire n_343, n_345, n_346, n_348, n_350, n_351, n_353, n_355;
  wire n_356, n_358, n_360, n_361, n_363, n_365, n_366, n_368;
  wire n_370, n_371, n_373, n_375, n_376, n_378, n_380, n_381;
  wire n_383, n_385, n_386, n_388, n_390, n_391, n_393, n_417;
  wire n_419, n_420, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445;
  and g1 (Z[0], A[0], B[0]);
  and g2 (n_46, A[1], B[0]);
  and g3 (n_63, A[2], B[0]);
  and g4 (n_67, A[3], B[0]);
  and g5 (n_72, A[4], B[0]);
  and g6 (n_80, A[5], B[0]);
  and g7 (n_90, A[6], B[0]);
  and g8 (n_103, A[7], B[0]);
  and g9 (n_61, A[0], B[1]);
  and g10 (n_45, A[1], B[1]);
  and g11 (n_68, A[2], B[1]);
  and g12 (n_73, A[3], B[1]);
  and g13 (n_64, A[4], B[1]);
  and g14 (n_91, A[5], B[1]);
  and g15 (n_104, A[6], B[1]);
  and g16 (n_120, A[7], B[1]);
  and g17 (n_66, A[0], B[2]);
  and g18 (n_70, A[1], B[2]);
  and g19 (n_76, A[2], B[2]);
  and g20 (n_83, A[3], B[2]);
  and g21 (n_94, A[4], B[2]);
  and g22 (n_108, A[5], B[2]);
  and g23 (n_121, A[6], B[2]);
  and g24 (n_137, A[7], B[2]);
  and g25 (n_69, A[0], B[3]);
  and g26 (n_74, A[1], B[3]);
  and g27 (n_81, A[2], B[3]);
  and g28 (n_92, A[3], B[3]);
  and g29 (n_105, A[4], B[3]);
  and g30 (n_124, A[5], B[3]);
  and g31 (n_138, A[6], B[3]);
  and g32 (n_152, A[7], B[3]);
  and g33 (n_75, A[0], B[4]);
  and g34 (n_82, A[1], B[4]);
  and g35 (n_93, A[2], B[4]);
  and g36 (n_107, A[3], B[4]);
  and g37 (n_122, A[4], B[4]);
  and g38 (n_141, A[5], B[4]);
  and g39 (n_153, A[6], B[4]);
  and g40 (n_164, A[7], B[4]);
  and g41 (n_84, A[0], B[5]);
  and g42 (n_65, A[1], B[5]);
  and g43 (n_109, A[2], B[5]);
  and g44 (n_123, A[3], B[5]);
  and g45 (n_139, A[4], B[5]);
  and g46 (n_156, A[5], B[5]);
  and g47 (n_165, A[6], B[5]);
  and g48 (n_173, A[7], B[5]);
  and g49 (n_95, A[0], B[6]);
  and g50 (n_110, A[1], B[6]);
  and g51 (n_125, A[2], B[6]);
  and g52 (n_140, A[3], B[6]);
  and g53 (n_154, A[4], B[6]);
  and g54 (n_167, A[5], B[6]);
  and g55 (n_174, A[6], B[6]);
  and g56 (n_179, A[7], B[6]);
  and g57 (n_106, A[0], B[7]);
  and g58 (n_126, A[1], B[7]);
  and g59 (n_142, A[2], B[7]);
  and g60 (n_155, A[3], B[7]);
  and g61 (n_166, A[4], B[7]);
  and g62 (n_175, A[5], B[7]);
  and g63 (n_180, A[6], B[7]);
  and g64 (n_33, A[7], B[7]);
  xor g107 (n_60, n_63, n_66);
  and g108 (n_44, n_63, n_66);
  xor g109 (n_71, n_67, n_68);
  and g110 (n_78, n_67, n_68);
  xor g111 (n_182, n_69, n_70);
  xor g112 (n_59, n_182, n_71);
  nand g113 (n_183, n_69, n_70);
  nand g114 (n_184, n_71, n_70);
  nand g115 (n_185, n_69, n_71);
  nand g116 (n_43, n_183, n_184, n_185);
  xor g117 (n_77, n_72, n_73);
  and g118 (n_86, n_72, n_73);
  xor g119 (n_186, n_74, n_75);
  xor g120 (n_79, n_186, n_76);
  nand g121 (n_187, n_74, n_75);
  nand g122 (n_188, n_76, n_75);
  nand g123 (n_189, n_74, n_76);
  nand g124 (n_87, n_187, n_188, n_189);
  xor g125 (n_190, n_77, n_78);
  xor g126 (n_58, n_190, n_79);
  nand g127 (n_191, n_77, n_78);
  nand g128 (n_192, n_79, n_78);
  nand g129 (n_193, n_77, n_79);
  nand g130 (n_42, n_191, n_192, n_193);
  xor g131 (n_85, n_80, n_64);
  and g132 (n_96, n_80, n_64);
  xor g133 (n_194, n_81, n_82);
  xor g134 (n_88, n_194, n_83);
  nand g135 (n_195, n_81, n_82);
  nand g136 (n_196, n_83, n_82);
  nand g137 (n_197, n_81, n_83);
  nand g138 (n_98, n_195, n_196, n_197);
  xor g139 (n_198, n_84, n_85);
  xor g140 (n_89, n_198, n_86);
  nand g141 (n_199, n_84, n_85);
  nand g142 (n_200, n_86, n_85);
  nand g143 (n_201, n_84, n_86);
  nand g144 (n_100, n_199, n_200, n_201);
  xor g145 (n_202, n_87, n_88);
  xor g146 (n_57, n_202, n_89);
  nand g147 (n_203, n_87, n_88);
  nand g148 (n_204, n_89, n_88);
  nand g149 (n_205, n_87, n_89);
  nand g150 (n_41, n_203, n_204, n_205);
  xor g151 (n_97, n_90, n_91);
  and g152 (n_111, n_90, n_91);
  xor g153 (n_206, n_92, n_93);
  xor g154 (n_99, n_206, n_94);
  nand g155 (n_207, n_92, n_93);
  nand g156 (n_208, n_94, n_93);
  nand g157 (n_209, n_92, n_94);
  nand g158 (n_113, n_207, n_208, n_209);
  xor g159 (n_210, n_65, n_95);
  xor g160 (n_101, n_210, n_96);
  nand g161 (n_211, n_65, n_95);
  nand g162 (n_212, n_96, n_95);
  nand g163 (n_213, n_65, n_96);
  nand g164 (n_116, n_211, n_212, n_213);
  xor g165 (n_214, n_97, n_98);
  xor g166 (n_102, n_214, n_99);
  nand g167 (n_215, n_97, n_98);
  nand g168 (n_216, n_99, n_98);
  nand g169 (n_217, n_97, n_99);
  nand g170 (n_118, n_215, n_216, n_217);
  xor g171 (n_218, n_100, n_101);
  xor g172 (n_56, n_218, n_102);
  nand g173 (n_219, n_100, n_101);
  nand g174 (n_220, n_102, n_101);
  nand g175 (n_221, n_100, n_102);
  nand g176 (n_40, n_219, n_220, n_221);
  xor g177 (n_112, n_103, n_104);
  and g178 (n_128, n_103, n_104);
  xor g179 (n_222, n_105, n_106);
  xor g180 (n_115, n_222, n_107);
  nand g181 (n_223, n_105, n_106);
  nand g182 (n_224, n_107, n_106);
  nand g183 (n_225, n_105, n_107);
  nand g184 (n_129, n_223, n_224, n_225);
  xor g185 (n_226, n_108, n_109);
  xor g186 (n_114, n_226, n_110);
  nand g187 (n_227, n_108, n_109);
  nand g188 (n_228, n_110, n_109);
  nand g189 (n_229, n_108, n_110);
  nand g190 (n_130, n_227, n_228, n_229);
  xor g191 (n_230, n_111, n_112);
  xor g192 (n_117, n_230, n_113);
  nand g193 (n_231, n_111, n_112);
  nand g194 (n_232, n_113, n_112);
  nand g195 (n_233, n_111, n_113);
  nand g196 (n_133, n_231, n_232, n_233);
  xor g197 (n_234, n_114, n_115);
  xor g198 (n_119, n_234, n_116);
  nand g199 (n_235, n_114, n_115);
  nand g200 (n_236, n_116, n_115);
  nand g201 (n_237, n_114, n_116);
  nand g202 (n_135, n_235, n_236, n_237);
  xor g203 (n_238, n_117, n_118);
  xor g204 (n_55, n_238, n_119);
  nand g205 (n_239, n_117, n_118);
  nand g206 (n_240, n_119, n_118);
  nand g207 (n_241, n_117, n_119);
  nand g208 (n_39, n_239, n_240, n_241);
  xor g209 (n_127, n_120, n_121);
  and g210 (n_143, n_120, n_121);
  xor g211 (n_242, n_122, n_123);
  xor g212 (n_131, n_242, n_124);
  nand g213 (n_243, n_122, n_123);
  nand g214 (n_244, n_124, n_123);
  nand g215 (n_245, n_122, n_124);
  nand g216 (n_144, n_243, n_244, n_245);
  xor g217 (n_246, n_125, n_126);
  xor g218 (n_132, n_246, n_127);
  nand g219 (n_247, n_125, n_126);
  nand g220 (n_248, n_127, n_126);
  nand g221 (n_249, n_125, n_127);
  nand g222 (n_147, n_247, n_248, n_249);
  xor g223 (n_250, n_128, n_129);
  xor g224 (n_134, n_250, n_130);
  nand g225 (n_251, n_128, n_129);
  nand g226 (n_252, n_130, n_129);
  nand g227 (n_253, n_128, n_130);
  nand g228 (n_148, n_251, n_252, n_253);
  xor g229 (n_254, n_131, n_132);
  xor g230 (n_136, n_254, n_133);
  nand g231 (n_255, n_131, n_132);
  nand g232 (n_256, n_133, n_132);
  nand g233 (n_257, n_131, n_133);
  nand g234 (n_151, n_255, n_256, n_257);
  xor g235 (n_258, n_134, n_135);
  xor g236 (n_54, n_258, n_136);
  nand g237 (n_259, n_134, n_135);
  nand g238 (n_260, n_136, n_135);
  nand g239 (n_261, n_134, n_136);
  nand g240 (n_38, n_259, n_260, n_261);
  xor g241 (n_262, n_137, n_138);
  xor g242 (n_146, n_262, n_139);
  nand g243 (n_263, n_137, n_138);
  nand g244 (n_264, n_139, n_138);
  nand g245 (n_265, n_137, n_139);
  nand g246 (n_158, n_263, n_264, n_265);
  xor g247 (n_266, n_140, n_141);
  xor g248 (n_145, n_266, n_142);
  nand g249 (n_267, n_140, n_141);
  nand g250 (n_268, n_142, n_141);
  nand g251 (n_269, n_140, n_142);
  nand g252 (n_157, n_267, n_268, n_269);
  xor g253 (n_270, n_143, n_144);
  xor g254 (n_149, n_270, n_145);
  nand g255 (n_271, n_143, n_144);
  nand g256 (n_272, n_145, n_144);
  nand g257 (n_273, n_143, n_145);
  nand g258 (n_161, n_271, n_272, n_273);
  xor g259 (n_274, n_146, n_147);
  xor g260 (n_150, n_274, n_148);
  nand g261 (n_275, n_146, n_147);
  nand g262 (n_276, n_148, n_147);
  nand g263 (n_277, n_146, n_148);
  nand g264 (n_163, n_275, n_276, n_277);
  xor g265 (n_278, n_149, n_150);
  xor g266 (n_53, n_278, n_151);
  nand g267 (n_279, n_149, n_150);
  nand g268 (n_280, n_151, n_150);
  nand g269 (n_281, n_149, n_151);
  nand g270 (n_37, n_279, n_280, n_281);
  xor g271 (n_282, n_152, n_153);
  xor g272 (n_159, n_282, n_154);
  nand g273 (n_283, n_152, n_153);
  nand g274 (n_284, n_154, n_153);
  nand g275 (n_285, n_152, n_154);
  nand g276 (n_168, n_283, n_284, n_285);
  xor g277 (n_286, n_155, n_156);
  xor g278 (n_160, n_286, n_157);
  nand g279 (n_287, n_155, n_156);
  nand g280 (n_288, n_157, n_156);
  nand g281 (n_289, n_155, n_157);
  nand g282 (n_170, n_287, n_288, n_289);
  xor g283 (n_290, n_158, n_159);
  xor g284 (n_162, n_290, n_160);
  nand g285 (n_291, n_158, n_159);
  nand g286 (n_292, n_160, n_159);
  nand g287 (n_293, n_158, n_160);
  nand g288 (n_172, n_291, n_292, n_293);
  xor g289 (n_294, n_161, n_162);
  xor g290 (n_52, n_294, n_163);
  nand g291 (n_295, n_161, n_162);
  nand g292 (n_296, n_163, n_162);
  nand g293 (n_297, n_161, n_163);
  nand g294 (n_36, n_295, n_296, n_297);
  xor g295 (n_298, n_164, n_165);
  xor g296 (n_169, n_298, n_166);
  nand g297 (n_299, n_164, n_165);
  nand g298 (n_300, n_166, n_165);
  nand g299 (n_301, n_164, n_166);
  nand g300 (n_176, n_299, n_300, n_301);
  xor g301 (n_302, n_167, n_168);
  xor g302 (n_171, n_302, n_169);
  nand g303 (n_303, n_167, n_168);
  nand g304 (n_304, n_169, n_168);
  nand g305 (n_305, n_167, n_169);
  nand g306 (n_178, n_303, n_304, n_305);
  xor g307 (n_306, n_170, n_171);
  xor g308 (n_51, n_306, n_172);
  nand g309 (n_307, n_170, n_171);
  nand g310 (n_308, n_172, n_171);
  nand g311 (n_309, n_170, n_172);
  nand g312 (n_50, n_307, n_308, n_309);
  xor g313 (n_310, n_173, n_174);
  xor g314 (n_177, n_310, n_175);
  nand g315 (n_311, n_173, n_174);
  nand g316 (n_312, n_175, n_174);
  nand g317 (n_313, n_173, n_175);
  nand g318 (n_181, n_311, n_312, n_313);
  xor g319 (n_314, n_176, n_177);
  xor g320 (n_35, n_314, n_178);
  nand g321 (n_315, n_176, n_177);
  nand g322 (n_316, n_178, n_177);
  nand g323 (n_317, n_176, n_178);
  nand g324 (n_49, n_315, n_316, n_317);
  xor g325 (n_318, n_179, n_180);
  xor g326 (n_34, n_318, n_181);
  nand g327 (n_319, n_179, n_180);
  nand g328 (n_320, n_181, n_180);
  nand g329 (n_321, n_179, n_181);
  nand g330 (n_48, n_319, n_320, n_321);
  nor g336 (n_325, n_46, n_61);
  nand g337 (n_328, n_46, n_61);
  nor g338 (n_330, n_45, n_60);
  nand g339 (n_333, n_45, n_60);
  nor g340 (n_335, n_44, n_59);
  nand g341 (n_338, n_44, n_59);
  nor g342 (n_340, n_43, n_58);
  nand g343 (n_343, n_43, n_58);
  nor g344 (n_345, n_42, n_57);
  nand g345 (n_348, n_42, n_57);
  nor g346 (n_350, n_41, n_56);
  nand g347 (n_353, n_41, n_56);
  nor g348 (n_355, n_40, n_55);
  nand g349 (n_358, n_40, n_55);
  nor g350 (n_360, n_39, n_54);
  nand g351 (n_363, n_39, n_54);
  nor g352 (n_365, n_38, n_53);
  nand g353 (n_368, n_38, n_53);
  nor g354 (n_370, n_37, n_52);
  nand g355 (n_373, n_37, n_52);
  nor g356 (n_375, n_36, n_51);
  nand g357 (n_378, n_36, n_51);
  nor g358 (n_380, n_35, n_50);
  nand g359 (n_383, n_35, n_50);
  nor g360 (n_385, n_34, n_49);
  nand g361 (n_388, n_34, n_49);
  nor g362 (n_390, n_33, n_48);
  nand g363 (n_393, n_33, n_48);
  nand g371 (n_336, n_333, n_420);
  nand g374 (n_341, n_338, n_424);
  nand g377 (n_346, n_343, n_428);
  nand g380 (n_351, n_348, n_434);
  nand g383 (n_356, n_353, n_437);
  nand g386 (n_361, n_358, n_438);
  nand g389 (n_366, n_363, n_439);
  nand g392 (n_371, n_368, n_440);
  nand g65 (n_376, n_373, n_441);
  nand g68 (n_381, n_378, n_442);
  nand g71 (n_386, n_383, n_443);
  nand g74 (n_391, n_388, n_444);
  nand g77 (Z[15], n_393, n_445);
  xnor g86 (Z[3], n_336, n_422);
  xnor g88 (Z[4], n_341, n_423);
  xnor g90 (Z[5], n_346, n_425);
  xnor g92 (Z[6], n_351, n_427);
  xnor g94 (Z[7], n_356, n_429);
  xnor g96 (Z[8], n_361, n_431);
  xnor g98 (Z[9], n_366, n_432);
  xnor g100 (Z[10], n_371, n_435);
  xnor g102 (Z[11], n_376, n_436);
  xnor g104 (Z[12], n_381, n_433);
  xnor g106 (Z[13], n_386, n_430);
  xnor g396 (Z[14], n_391, n_426);
  or g400 (n_417, wc, n_325);
  not gc (wc, n_328);
  not g402 (Z[1], n_417);
  or g403 (n_419, wc0, n_330);
  not gc0 (wc0, n_333);
  or g404 (n_420, n_328, n_330);
  xor g405 (Z[2], n_328, n_419);
  or g406 (n_422, wc1, n_335);
  not gc1 (wc1, n_338);
  or g407 (n_423, wc2, n_340);
  not gc2 (wc2, n_343);
  or g408 (n_424, wc3, n_335);
  not gc3 (wc3, n_336);
  or g409 (n_425, wc4, n_345);
  not gc4 (wc4, n_348);
  or g410 (n_426, wc5, n_390);
  not gc5 (wc5, n_393);
  or g411 (n_427, wc6, n_350);
  not gc6 (wc6, n_353);
  or g412 (n_428, wc7, n_340);
  not gc7 (wc7, n_341);
  or g413 (n_429, wc8, n_355);
  not gc8 (wc8, n_358);
  or g414 (n_430, wc9, n_385);
  not gc9 (wc9, n_388);
  or g415 (n_431, wc10, n_360);
  not gc10 (wc10, n_363);
  or g416 (n_432, wc11, n_365);
  not gc11 (wc11, n_368);
  or g417 (n_433, wc12, n_380);
  not gc12 (wc12, n_383);
  or g418 (n_434, wc13, n_345);
  not gc13 (wc13, n_346);
  or g419 (n_435, wc14, n_370);
  not gc14 (wc14, n_373);
  or g420 (n_436, wc15, n_375);
  not gc15 (wc15, n_378);
  or g421 (n_437, wc16, n_350);
  not gc16 (wc16, n_351);
  or g422 (n_438, wc17, n_355);
  not gc17 (wc17, n_356);
  or g423 (n_439, wc18, n_360);
  not gc18 (wc18, n_361);
  or g424 (n_440, wc19, n_365);
  not gc19 (wc19, n_366);
  or g425 (n_441, wc20, n_370);
  not gc20 (wc20, n_371);
  or g426 (n_442, wc21, n_375);
  not gc21 (wc21, n_376);
  or g427 (n_443, wc22, n_380);
  not gc22 (wc22, n_381);
  or g428 (n_444, wc23, n_385);
  not gc23 (wc23, n_386);
  or g429 (n_445, wc24, n_390);
  not gc24 (wc24, n_391);
endmodule

module mult_unsigned_GENERIC(A, B, Z);
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  mult_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

