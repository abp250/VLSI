library verilog;
use verilog.vl_types.all;
entity Elevator_tb is
end Elevator_tb;
