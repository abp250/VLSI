library verilog;
use verilog.vl_types.all;
entity t_control is
end t_control;
