module add_unsigned_carry_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_unsigned_carry
  input [16:0] A, B;
  input CI;
  output [16:0] Z;
  wire [16:0] A, B;
  wire CI;
  wire [16:0] Z;
  wire n_53, n_54, n_55, n_56, n_57, n_59, n_61, n_62;
  wire n_63, n_64, n_66, n_67, n_68, n_69, n_70, n_72;
  wire n_73, n_74, n_75, n_76, n_78, n_79, n_80, n_81;
  wire n_82, n_84, n_85, n_86, n_87, n_88, n_90, n_91;
  wire n_92, n_93, n_94, n_96, n_97, n_98, n_99, n_100;
  wire n_102, n_103, n_106, n_108, n_109, n_110, n_112, n_114;
  wire n_119, n_120, n_122, n_124, n_129, n_130, n_132, n_134;
  wire n_139, n_142, n_147, n_151, n_152, n_154, n_158, n_160;
  wire n_162, n_164, n_166, n_169, n_176, n_178, n_181, n_182;
  wire n_184, n_185, n_187, n_188, n_189, n_191, n_196, n_200;
  wire n_202, n_205, n_209, n_211, n_214, n_217, n_220, n_222;
  wire n_225, n_228, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277;
  xor g1 (n_228, A[0], B[0]);
  nand g2 (n_53, A[0], B[0]);
  nand g3 (n_54, A[0], CI);
  nand g4 (n_55, B[0], CI);
  nand g5 (n_57, n_53, n_54, n_55);
  nor g6 (n_56, A[1], B[1]);
  nand g7 (n_59, A[1], B[1]);
  nor g8 (n_66, A[2], B[2]);
  nand g9 (n_61, A[2], B[2]);
  nor g10 (n_62, A[3], B[3]);
  nand g11 (n_63, A[3], B[3]);
  nor g12 (n_72, A[4], B[4]);
  nand g13 (n_67, A[4], B[4]);
  nor g14 (n_68, A[5], B[5]);
  nand g15 (n_69, A[5], B[5]);
  nor g16 (n_78, A[6], B[6]);
  nand g17 (n_73, A[6], B[6]);
  nor g18 (n_74, A[7], B[7]);
  nand g19 (n_75, A[7], B[7]);
  nor g20 (n_84, A[8], B[8]);
  nand g21 (n_79, A[8], B[8]);
  nor g22 (n_80, A[9], B[9]);
  nand g23 (n_81, A[9], B[9]);
  nor g24 (n_90, A[10], B[10]);
  nand g25 (n_85, A[10], B[10]);
  nor g26 (n_86, A[11], B[11]);
  nand g27 (n_87, A[11], B[11]);
  nor g28 (n_96, A[12], B[12]);
  nand g29 (n_91, A[12], B[12]);
  nor g30 (n_92, A[13], B[13]);
  nand g31 (n_93, A[13], B[13]);
  nor g32 (n_102, A[14], B[14]);
  nand g33 (n_97, A[14], B[14]);
  nor g34 (n_98, A[15], B[15]);
  nand g35 (n_99, A[15], B[15]);
  nor g36 (n_188, A[16], B[16]);
  nand g37 (n_191, A[16], B[16]);
  nand g40 (n_103, n_59, n_234);
  nor g41 (n_64, n_61, n_62);
  nor g44 (n_106, n_66, n_62);
  nor g45 (n_70, n_67, n_68);
  nor g48 (n_112, n_72, n_68);
  nor g49 (n_76, n_73, n_74);
  nor g52 (n_114, n_78, n_74);
  nor g53 (n_82, n_79, n_80);
  nor g56 (n_122, n_84, n_80);
  nor g57 (n_88, n_85, n_86);
  nor g60 (n_124, n_90, n_86);
  nor g61 (n_94, n_91, n_92);
  nor g64 (n_132, n_96, n_92);
  nor g65 (n_100, n_97, n_98);
  nor g68 (n_134, n_102, n_98);
  nand g71 (n_196, n_61, n_261);
  nand g72 (n_108, n_106, n_103);
  nand g73 (n_139, n_235, n_108);
  nor g74 (n_110, n_78, n_109);
  nand g83 (n_147, n_112, n_114);
  nor g84 (n_120, n_90, n_119);
  nand g93 (n_154, n_122, n_124);
  nor g94 (n_130, n_102, n_129);
  nand g103 (n_162, n_132, n_134);
  nand g106 (n_200, n_67, n_268);
  nand g107 (n_142, n_112, n_139);
  nand g108 (n_202, n_109, n_142);
  nand g111 (n_205, n_262, n_269);
  nand g114 (n_166, n_263, n_270);
  nor g115 (n_152, n_96, n_151);
  nor g118 (n_176, n_96, n_154);
  nor g124 (n_160, n_158, n_151);
  nor g127 (n_182, n_154, n_158);
  nor g128 (n_164, n_162, n_151);
  nor g131 (n_185, n_154, n_162);
  nand g134 (n_209, n_79, n_275);
  nand g135 (n_169, n_122, n_166);
  nand g136 (n_211, n_119, n_169);
  nand g139 (n_214, n_264, n_276);
  nand g142 (n_217, n_151, n_277);
  nand g143 (n_178, n_176, n_166);
  nand g144 (n_220, n_271, n_178);
  nand g145 (n_181, n_260, n_166);
  nand g146 (n_222, n_272, n_181);
  nand g147 (n_184, n_182, n_166);
  nand g148 (n_225, n_273, n_184);
  nand g149 (n_187, n_185, n_166);
  nand g150 (n_189, n_274, n_187);
  xnor g155 (Z[1], n_57, n_241);
  xnor g157 (Z[2], n_103, n_242);
  xnor g160 (Z[3], n_196, n_243);
  xnor g162 (Z[4], n_139, n_244);
  xnor g165 (Z[5], n_200, n_245);
  xnor g167 (Z[6], n_202, n_246);
  xnor g170 (Z[7], n_205, n_247);
  xnor g172 (Z[8], n_166, n_248);
  xnor g175 (Z[9], n_209, n_249);
  xnor g177 (Z[10], n_211, n_250);
  xnor g180 (Z[11], n_214, n_251);
  xnor g183 (Z[12], n_217, n_252);
  xnor g186 (Z[13], n_220, n_253);
  xnor g188 (Z[14], n_222, n_254);
  xnor g191 (Z[15], n_225, n_255);
  xnor g193 (Z[16], n_189, n_256);
  xor g194 (Z[0], CI, n_228);
  or g195 (n_234, n_56, wc);
  not gc (wc, n_57);
  and g196 (n_235, wc0, n_63);
  not gc0 (wc0, n_64);
  and g197 (n_109, wc1, n_69);
  not gc1 (wc1, n_70);
  and g198 (n_236, wc2, n_75);
  not gc2 (wc2, n_76);
  and g199 (n_119, wc3, n_81);
  not gc3 (wc3, n_82);
  and g200 (n_237, wc4, n_87);
  not gc4 (wc4, n_88);
  and g201 (n_129, wc5, n_93);
  not gc5 (wc5, n_94);
  and g202 (n_238, wc6, n_99);
  not gc6 (wc6, n_100);
  or g203 (n_239, wc7, n_78);
  not gc7 (wc7, n_112);
  or g204 (n_240, wc8, n_90);
  not gc8 (wc8, n_122);
  or g205 (n_158, wc9, n_102);
  not gc9 (wc9, n_132);
  or g206 (n_241, wc10, n_56);
  not gc10 (wc10, n_59);
  or g207 (n_242, wc11, n_66);
  not gc11 (wc11, n_61);
  or g208 (n_243, wc12, n_62);
  not gc12 (wc12, n_63);
  or g209 (n_244, wc13, n_72);
  not gc13 (wc13, n_67);
  or g210 (n_245, wc14, n_68);
  not gc14 (wc14, n_69);
  or g211 (n_246, wc15, n_78);
  not gc15 (wc15, n_73);
  or g212 (n_247, wc16, n_74);
  not gc16 (wc16, n_75);
  or g213 (n_248, wc17, n_84);
  not gc17 (wc17, n_79);
  or g214 (n_249, wc18, n_80);
  not gc18 (wc18, n_81);
  or g215 (n_250, wc19, n_90);
  not gc19 (wc19, n_85);
  or g216 (n_251, wc20, n_86);
  not gc20 (wc20, n_87);
  or g217 (n_252, wc21, n_96);
  not gc21 (wc21, n_91);
  or g218 (n_253, wc22, n_92);
  not gc22 (wc22, n_93);
  or g219 (n_254, wc23, n_102);
  not gc23 (wc23, n_97);
  or g220 (n_255, wc24, n_98);
  not gc24 (wc24, n_99);
  or g221 (n_256, wc25, n_188);
  not gc25 (wc25, n_191);
  and g222 (n_257, wc26, n_114);
  not gc26 (wc26, n_109);
  and g223 (n_258, wc27, n_124);
  not gc27 (wc27, n_119);
  and g224 (n_259, wc28, n_134);
  not gc28 (wc28, n_129);
  and g225 (n_260, wc29, n_132);
  not gc29 (wc29, n_154);
  or g226 (n_261, wc30, n_66);
  not gc30 (wc30, n_103);
  and g227 (n_262, wc31, n_73);
  not gc31 (wc31, n_110);
  and g228 (n_263, wc32, n_236);
  not gc32 (wc32, n_257);
  and g229 (n_264, wc33, n_85);
  not gc33 (wc33, n_120);
  and g230 (n_151, wc34, n_237);
  not gc34 (wc34, n_258);
  and g231 (n_265, wc35, n_97);
  not gc35 (wc35, n_130);
  and g232 (n_266, wc36, n_238);
  not gc36 (wc36, n_259);
  and g233 (n_267, wc37, n_132);
  not gc37 (wc37, n_151);
  or g234 (n_268, wc38, n_72);
  not gc38 (wc38, n_139);
  or g235 (n_269, n_239, wc39);
  not gc39 (wc39, n_139);
  or g236 (n_270, n_147, wc40);
  not gc40 (wc40, n_139);
  and g237 (n_271, wc41, n_91);
  not gc41 (wc41, n_152);
  and g238 (n_272, wc42, n_129);
  not gc42 (wc42, n_267);
  and g239 (n_273, n_265, wc43);
  not gc43 (wc43, n_160);
  and g240 (n_274, n_266, wc44);
  not gc44 (wc44, n_164);
  or g241 (n_275, wc45, n_84);
  not gc45 (wc45, n_166);
  or g242 (n_276, n_240, wc46);
  not gc46 (wc46, n_166);
  or g243 (n_277, wc47, n_154);
  not gc47 (wc47, n_166);
endmodule

module add_unsigned_carry_GENERIC(A, B, CI, Z);
  input [16:0] A, B;
  input CI;
  output [16:0] Z;
  wire [16:0] A, B;
  wire CI;
  wire [16:0] Z;
  add_unsigned_carry_GENERIC_REAL g1(.A (A), .B (B), .CI (CI), .Z (Z));
endmodule

module bmux_1_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [16:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  or g18 (z[16], wc, wc1);
  and gc1 (wc1, in_1[16], ctl);
  and gc0 (wc, in_0[16], wc0);
  not gc (wc0, ctl);
  or g19 (z[15], wc2, wc4);
  and gc4 (wc4, in_1[15], ctl);
  and gc3 (wc2, in_0[15], wc3);
  not gc2 (wc3, ctl);
  or g20 (z[14], wc5, wc7);
  and gc7 (wc7, in_1[14], ctl);
  and gc6 (wc5, in_0[14], wc6);
  not gc5 (wc6, ctl);
  or g21 (z[13], wc8, wc10);
  and gc10 (wc10, in_1[13], ctl);
  and gc9 (wc8, in_0[13], wc9);
  not gc8 (wc9, ctl);
  or g22 (z[12], wc11, wc13);
  and gc13 (wc13, in_1[12], ctl);
  and gc12 (wc11, in_0[12], wc12);
  not gc11 (wc12, ctl);
  or g23 (z[11], wc14, wc16);
  and gc16 (wc16, in_1[11], ctl);
  and gc15 (wc14, in_0[11], wc15);
  not gc14 (wc15, ctl);
  or g24 (z[10], wc17, wc19);
  and gc19 (wc19, in_1[10], ctl);
  and gc18 (wc17, in_0[10], wc18);
  not gc17 (wc18, ctl);
  or g25 (z[9], wc20, wc22);
  and gc22 (wc22, in_1[9], ctl);
  and gc21 (wc20, in_0[9], wc21);
  not gc20 (wc21, ctl);
  or g26 (z[8], wc23, wc25);
  and gc25 (wc25, in_1[8], ctl);
  and gc24 (wc23, in_0[8], wc24);
  not gc23 (wc24, ctl);
  or g27 (z[7], wc26, wc28);
  and gc28 (wc28, in_1[7], ctl);
  and gc27 (wc26, in_0[7], wc27);
  not gc26 (wc27, ctl);
  or g28 (z[6], wc29, wc31);
  and gc31 (wc31, in_1[6], ctl);
  and gc30 (wc29, in_0[6], wc30);
  not gc29 (wc30, ctl);
  or g29 (z[5], wc32, wc34);
  and gc34 (wc34, in_1[5], ctl);
  and gc33 (wc32, in_0[5], wc33);
  not gc32 (wc33, ctl);
  or g30 (z[4], wc35, wc37);
  and gc37 (wc37, in_1[4], ctl);
  and gc36 (wc35, in_0[4], wc36);
  not gc35 (wc36, ctl);
  or g31 (z[3], wc38, wc40);
  and gc40 (wc40, in_1[3], ctl);
  and gc39 (wc38, in_0[3], wc39);
  not gc38 (wc39, ctl);
  or g32 (z[2], wc41, wc43);
  and gc43 (wc43, in_1[2], ctl);
  and gc42 (wc41, in_0[2], wc42);
  not gc41 (wc42, ctl);
  or g33 (z[1], wc44, wc46);
  and gc46 (wc46, in_1[1], ctl);
  and gc45 (wc44, in_0[1], wc45);
  not gc44 (wc45, ctl);
  or g34 (z[0], wc47, wc49);
  and gc49 (wc49, in_1[0], ctl);
  and gc48 (wc47, in_0[0], wc48);
  not gc47 (wc48, ctl);
endmodule

module bmux_1_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  bmux_1_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1), .z
       (z));
endmodule

module bmux_2_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [16:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  or g18 (z[16], wc, wc1);
  and gc1 (wc1, in_1[16], ctl);
  and gc0 (wc, in_0[16], wc0);
  not gc (wc0, ctl);
  or g19 (z[15], wc2, wc4);
  and gc4 (wc4, in_1[15], ctl);
  and gc3 (wc2, in_0[15], wc3);
  not gc2 (wc3, ctl);
  or g20 (z[14], wc5, wc7);
  and gc7 (wc7, in_1[14], ctl);
  and gc6 (wc5, in_0[14], wc6);
  not gc5 (wc6, ctl);
  or g21 (z[13], wc8, wc10);
  and gc10 (wc10, in_1[13], ctl);
  and gc9 (wc8, in_0[13], wc9);
  not gc8 (wc9, ctl);
  or g22 (z[12], wc11, wc13);
  and gc13 (wc13, in_1[12], ctl);
  and gc12 (wc11, in_0[12], wc12);
  not gc11 (wc12, ctl);
  or g23 (z[11], wc14, wc16);
  and gc16 (wc16, in_1[11], ctl);
  and gc15 (wc14, in_0[11], wc15);
  not gc14 (wc15, ctl);
  or g24 (z[10], wc17, wc19);
  and gc19 (wc19, in_1[10], ctl);
  and gc18 (wc17, in_0[10], wc18);
  not gc17 (wc18, ctl);
  or g25 (z[9], wc20, wc22);
  and gc22 (wc22, in_1[9], ctl);
  and gc21 (wc20, in_0[9], wc21);
  not gc20 (wc21, ctl);
  or g26 (z[8], wc23, wc25);
  and gc25 (wc25, in_1[8], ctl);
  and gc24 (wc23, in_0[8], wc24);
  not gc23 (wc24, ctl);
  or g27 (z[7], wc26, wc28);
  and gc28 (wc28, in_1[7], ctl);
  and gc27 (wc26, in_0[7], wc27);
  not gc26 (wc27, ctl);
  or g28 (z[6], wc29, wc31);
  and gc31 (wc31, in_1[6], ctl);
  and gc30 (wc29, in_0[6], wc30);
  not gc29 (wc30, ctl);
  or g29 (z[5], wc32, wc34);
  and gc34 (wc34, in_1[5], ctl);
  and gc33 (wc32, in_0[5], wc33);
  not gc32 (wc33, ctl);
  or g30 (z[4], wc35, wc37);
  and gc37 (wc37, in_1[4], ctl);
  and gc36 (wc35, in_0[4], wc36);
  not gc35 (wc36, ctl);
  or g31 (z[3], wc38, wc40);
  and gc40 (wc40, in_1[3], ctl);
  and gc39 (wc38, in_0[3], wc39);
  not gc38 (wc39, ctl);
  or g32 (z[2], wc41, wc43);
  and gc43 (wc43, in_1[2], ctl);
  and gc42 (wc41, in_0[2], wc42);
  not gc41 (wc42, ctl);
  or g33 (z[1], wc44, wc46);
  and gc46 (wc46, in_1[1], ctl);
  and gc45 (wc44, in_0[1], wc45);
  not gc44 (wc45, ctl);
  or g34 (z[0], wc47, wc49);
  and gc49 (wc49, in_1[0], ctl);
  and gc48 (wc47, in_0[0], wc48);
  not gc47 (wc48, ctl);
endmodule

module bmux_2_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [16:0] in_0, in_1;
  output [16:0] z;
  wire ctl;
  wire [16:0] in_0, in_1;
  wire [16:0] z;
  bmux_2_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1), .z
       (z));
endmodule

module bmux_50_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [0:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl, in_0, in_1;
  output z;
  wire ctl, in_0, in_1;
  wire z;
  or g2 (z, wc, wc1);
  and gc1 (wc1, in_1, ctl);
  and gc0 (wc, in_0, wc0);
  not gc (wc0, ctl);
endmodule

module bmux_50_GENERIC(ctl, in_0, in_1, z);
  input ctl, in_0, in_1;
  output z;
  wire ctl, in_0, in_1;
  wire z;
  bmux_50_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1), .z
       (z));
endmodule

module csa_tree_GENERIC_REAL(in_0, in_1, in_2, in_3, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( in_0 * in_1 )  + ( in_2 * in_3 )  )  ; assign out_1 = 17'b0;"
  input [7:0] in_0, in_1, in_2, in_3;
  output [16:0] out_0, out_1;
  wire [7:0] in_0, in_1, in_2, in_3;
  wire [16:0] out_0, out_1;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697;
  wire n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  assign out_1[16] = 1'b0;
  assign out_0[16] = 1'b0;
  and g1 (out_0[0], in_0[0], in_1[0]);
  and g2 (n_33, in_0[1], in_1[0]);
  and g3 (n_36, in_0[2], in_1[0]);
  and g4 (n_44, in_0[3], in_1[0]);
  and g5 (n_58, in_0[4], in_1[0]);
  and g6 (n_78, in_0[5], in_1[0]);
  and g7 (n_104, in_0[6], in_1[0]);
  and g8 (n_136, in_0[7], in_1[0]);
  and g9 (out_0[1], in_0[0], in_1[1]);
  and g10 (n_37, in_0[1], in_1[1]);
  and g11 (n_45, in_0[2], in_1[1]);
  and g12 (n_59, in_0[3], in_1[1]);
  and g13 (n_79, in_0[4], in_1[1]);
  and g14 (n_105, in_0[5], in_1[1]);
  and g15 (n_137, in_0[6], in_1[1]);
  and g16 (n_174, in_0[7], in_1[1]);
  and g17 (n_41, in_0[0], in_1[2]);
  and g18 (n_49, in_0[1], in_1[2]);
  and g19 (n_65, in_0[2], in_1[2]);
  and g20 (n_86, in_0[3], in_1[2]);
  and g21 (n_112, in_0[4], in_1[2]);
  and g22 (n_145, in_0[5], in_1[2]);
  and g23 (n_175, in_0[6], in_1[2]);
  and g24 (n_212, in_0[7], in_1[2]);
  and g25 (n_46, in_0[0], in_1[3]);
  and g26 (n_60, in_0[1], in_1[3]);
  and g27 (n_80, in_0[2], in_1[3]);
  and g28 (n_106, in_0[3], in_1[3]);
  and g29 (n_138, in_0[4], in_1[3]);
  and g30 (n_182, in_0[5], in_1[3]);
  and g31 (n_213, in_0[6], in_1[3]);
  and g32 (n_247, in_0[7], in_1[3]);
  and g33 (n_63, in_0[0], in_1[4]);
  and g34 (n_83, in_0[1], in_1[4]);
  and g35 (n_109, in_0[2], in_1[4]);
  and g36 (n_142, in_0[3], in_1[4]);
  and g37 (n_176, in_0[4], in_1[4]);
  and g38 (n_220, in_0[5], in_1[4]);
  and g39 (n_248, in_0[6], in_1[4]);
  and g40 (n_277, in_0[7], in_1[4]);
  and g41 (n_87, in_0[0], in_1[5]);
  and g42 (n_113, in_0[1], in_1[5]);
  and g43 (n_146, in_0[2], in_1[5]);
  and g44 (n_179, in_0[3], in_1[5]);
  and g45 (n_214, in_0[4], in_1[5]);
  and g46 (n_254, in_0[5], in_1[5]);
  and g47 (n_278, in_0[6], in_1[5]);
  and g48 (n_301, in_0[7], in_1[5]);
  and g49 (n_116, in_0[0], in_1[6]);
  and g50 (n_149, in_0[1], in_1[6]);
  and g51 (n_183, in_0[2], in_1[6]);
  and g52 (n_217, in_0[3], in_1[6]);
  and g53 (n_249, in_0[4], in_1[6]);
  and g54 (n_282, in_0[5], in_1[6]);
  and g55 (n_302, in_0[6], in_1[6]);
  and g56 (n_319, in_0[7], in_1[6]);
  and g57 (n_139, in_0[0], in_1[7]);
  and g58 (n_186, in_0[1], in_1[7]);
  and g59 (n_221, in_0[2], in_1[7]);
  and g60 (n_252, in_0[3], in_1[7]);
  and g61 (n_279, in_0[4], in_1[7]);
  and g62 (n_305, in_0[5], in_1[7]);
  and g63 (n_320, in_0[6], in_1[7]);
  and g64 (n_331, in_0[7], in_1[7]);
  and g65 (out_1[0], in_2[0], in_3[0]);
  and g66 (n_35, in_2[1], in_3[0]);
  and g67 (n_39, in_2[2], in_3[0]);
  and g68 (n_48, in_2[3], in_3[0]);
  and g69 (n_66, in_2[4], in_3[0]);
  and g70 (n_89, in_2[5], in_3[0]);
  and g71 (n_107, in_2[6], in_3[0]);
  and g72 (n_141, in_2[7], in_3[0]);
  and g73 (n_34, in_2[0], in_3[1]);
  and g74 (n_40, in_2[1], in_3[1]);
  and g75 (n_50, in_2[2], in_3[1]);
  and g76 (n_67, in_2[3], in_3[1]);
  and g77 (n_81, in_2[4], in_3[1]);
  and g78 (n_108, in_2[5], in_3[1]);
  and g79 (n_143, in_2[6], in_3[1]);
  and g80 (n_177, in_2[7], in_3[1]);
  and g81 (n_38, in_2[0], in_3[2]);
  and g82 (n_51, in_2[1], in_3[2]);
  and g83 (n_61, in_2[2], in_3[2]);
  and g84 (n_82, in_2[3], in_3[2]);
  and g85 (n_110, in_2[4], in_3[2]);
  and g86 (n_144, in_2[5], in_3[2]);
  and g87 (n_178, in_2[6], in_3[2]);
  and g88 (n_223, in_2[7], in_3[2]);
  and g89 (n_47, in_2[0], in_3[3]);
  and g90 (n_62, in_2[1], in_3[3]);
  and g91 (n_84, in_2[2], in_3[3]);
  and g92 (n_111, in_2[3], in_3[3]);
  and g93 (n_147, in_2[4], in_3[3]);
  and g94 (n_180, in_2[5], in_3[3]);
  and g95 (n_215, in_2[6], in_3[3]);
  and g96 (n_255, in_2[7], in_3[3]);
  and g97 (n_64, in_2[0], in_3[4]);
  and g98 (n_85, in_2[1], in_3[4]);
  and g99 (n_114, in_2[2], in_3[4]);
  and g100 (n_148, in_2[3], in_3[4]);
  and g101 (n_181, in_2[4], in_3[4]);
  and g102 (n_216, in_2[5], in_3[4]);
  and g103 (n_256, in_2[6], in_3[4]);
  and g104 (n_281, in_2[7], in_3[4]);
  and g105 (n_88, in_2[0], in_3[5]);
  and g106 (n_115, in_2[1], in_3[5]);
  and g107 (n_150, in_2[2], in_3[5]);
  and g108 (n_184, in_2[3], in_3[5]);
  and g109 (n_218, in_2[4], in_3[5]);
  and g110 (n_250, in_2[5], in_3[5]);
  and g111 (n_283, in_2[6], in_3[5]);
  and g112 (n_303, in_2[7], in_3[5]);
  and g113 (n_117, in_2[0], in_3[6]);
  and g114 (n_151, in_2[1], in_3[6]);
  and g115 (n_185, in_2[2], in_3[6]);
  and g116 (n_219, in_2[3], in_3[6]);
  and g117 (n_251, in_2[4], in_3[6]);
  and g118 (n_284, in_2[5], in_3[6]);
  and g119 (n_304, in_2[6], in_3[6]);
  and g120 (n_322, in_2[7], in_3[6]);
  and g121 (n_140, in_2[0], in_3[7]);
  and g122 (n_187, in_2[1], in_3[7]);
  and g123 (n_222, in_2[2], in_3[7]);
  and g124 (n_253, in_2[3], in_3[7]);
  and g125 (n_280, in_2[4], in_3[7]);
  and g126 (n_306, in_2[5], in_3[7]);
  and g127 (n_321, in_2[6], in_3[7]);
  and g128 (n_332, in_2[7], in_3[7]);
  xor g233 (n_370, n_33, n_34);
  xor g234 (out_1[1], n_370, n_35);
  nand g235 (n_371, n_33, n_34);
  nand g236 (n_372, n_35, n_34);
  nand g237 (n_373, n_33, n_35);
  nand g238 (n_43, n_371, n_372, n_373);
  xor g239 (n_42, n_36, n_37);
  and g240 (n_52, n_36, n_37);
  xor g241 (n_374, n_38, n_39);
  xor g242 (out_0[2], n_374, n_40);
  nand g243 (n_375, n_38, n_39);
  nand g244 (n_376, n_40, n_39);
  nand g245 (n_377, n_38, n_40);
  nand g246 (n_54, n_375, n_376, n_377);
  xor g247 (n_378, n_41, n_42);
  xor g248 (out_1[2], n_378, n_43);
  nand g249 (n_379, n_41, n_42);
  nand g250 (n_380, n_43, n_42);
  nand g251 (n_381, n_41, n_43);
  nand g252 (out_0[3], n_379, n_380, n_381);
  xor g253 (n_53, n_44, n_45);
  and g254 (n_69, n_44, n_45);
  xor g255 (n_382, n_46, n_47);
  xor g256 (n_56, n_382, n_48);
  nand g257 (n_383, n_46, n_47);
  nand g258 (n_384, n_48, n_47);
  nand g259 (n_385, n_46, n_48);
  nand g260 (n_70, n_383, n_384, n_385);
  xor g261 (n_386, n_49, n_50);
  xor g262 (n_55, n_386, n_51);
  nand g263 (n_387, n_49, n_50);
  nand g264 (n_388, n_51, n_50);
  nand g265 (n_389, n_49, n_51);
  nand g266 (n_71, n_387, n_388, n_389);
  xor g267 (n_390, n_52, n_53);
  xor g268 (n_57, n_390, n_54);
  nand g269 (n_391, n_52, n_53);
  nand g270 (n_392, n_54, n_53);
  nand g271 (n_393, n_52, n_54);
  nand g272 (n_75, n_391, n_392, n_393);
  xor g273 (n_394, n_55, n_56);
  xor g274 (out_1[3], n_394, n_57);
  nand g275 (n_395, n_55, n_56);
  nand g276 (n_396, n_57, n_56);
  nand g277 (n_397, n_55, n_57);
  nand g278 (out_0[4], n_395, n_396, n_397);
  xor g279 (n_68, n_58, n_59);
  and g280 (n_91, n_58, n_59);
  xor g281 (n_398, n_60, n_61);
  xor g282 (n_72, n_398, n_62);
  nand g283 (n_399, n_60, n_61);
  nand g284 (n_400, n_62, n_61);
  nand g285 (n_401, n_60, n_62);
  nand g286 (n_93, n_399, n_400, n_401);
  xor g287 (n_402, n_63, n_64);
  xor g288 (n_73, n_402, n_65);
  nand g289 (n_403, n_63, n_64);
  nand g290 (n_404, n_65, n_64);
  nand g291 (n_405, n_63, n_65);
  nand g292 (n_92, n_403, n_404, n_405);
  xor g293 (n_406, n_66, n_67);
  xor g294 (n_74, n_406, n_68);
  nand g295 (n_407, n_66, n_67);
  nand g296 (n_408, n_68, n_67);
  nand g297 (n_409, n_66, n_68);
  nand g298 (n_97, n_407, n_408, n_409);
  xor g299 (n_410, n_69, n_70);
  xor g300 (n_76, n_410, n_71);
  nand g301 (n_411, n_69, n_70);
  nand g302 (n_412, n_71, n_70);
  nand g303 (n_413, n_69, n_71);
  nand g304 (n_98, n_411, n_412, n_413);
  xor g305 (n_414, n_72, n_73);
  xor g306 (n_77, n_414, n_74);
  nand g307 (n_415, n_72, n_73);
  nand g308 (n_416, n_74, n_73);
  nand g309 (n_417, n_72, n_74);
  nand g310 (n_101, n_415, n_416, n_417);
  xor g311 (n_418, n_75, n_76);
  xor g312 (out_1[4], n_418, n_77);
  nand g313 (n_419, n_75, n_76);
  nand g314 (n_420, n_77, n_76);
  nand g315 (n_421, n_75, n_77);
  nand g316 (out_0[5], n_419, n_420, n_421);
  xor g317 (n_90, n_78, n_79);
  and g318 (n_119, n_78, n_79);
  xor g319 (n_422, n_80, n_81);
  xor g320 (n_95, n_422, n_82);
  nand g321 (n_423, n_80, n_81);
  nand g322 (n_424, n_82, n_81);
  nand g323 (n_425, n_80, n_82);
  nand g324 (n_120, n_423, n_424, n_425);
  xor g325 (n_426, n_83, n_84);
  xor g326 (n_96, n_426, n_85);
  nand g327 (n_427, n_83, n_84);
  nand g328 (n_428, n_85, n_84);
  nand g329 (n_429, n_83, n_85);
  nand g330 (n_121, n_427, n_428, n_429);
  xor g331 (n_430, n_86, n_87);
  xor g332 (n_94, n_430, n_88);
  nand g333 (n_431, n_86, n_87);
  nand g334 (n_432, n_88, n_87);
  nand g335 (n_433, n_86, n_88);
  nand g336 (n_122, n_431, n_432, n_433);
  xor g337 (n_434, n_89, n_90);
  xor g338 (n_99, n_434, n_91);
  nand g339 (n_435, n_89, n_90);
  nand g340 (n_436, n_91, n_90);
  nand g341 (n_437, n_89, n_91);
  nand g342 (n_127, n_435, n_436, n_437);
  xor g343 (n_438, n_92, n_93);
  xor g344 (n_100, n_438, n_94);
  nand g345 (n_439, n_92, n_93);
  nand g346 (n_440, n_94, n_93);
  nand g347 (n_441, n_92, n_94);
  nand g348 (n_130, n_439, n_440, n_441);
  xor g349 (n_442, n_95, n_96);
  xor g350 (n_102, n_442, n_97);
  nand g351 (n_443, n_95, n_96);
  nand g352 (n_444, n_97, n_96);
  nand g353 (n_445, n_95, n_97);
  nand g354 (n_132, n_443, n_444, n_445);
  xor g355 (n_446, n_98, n_99);
  xor g356 (n_103, n_446, n_100);
  nand g357 (n_447, n_98, n_99);
  nand g358 (n_448, n_100, n_99);
  nand g359 (n_449, n_98, n_100);
  nand g360 (n_134, n_447, n_448, n_449);
  xor g361 (n_450, n_101, n_102);
  xor g362 (out_1[5], n_450, n_103);
  nand g363 (n_451, n_101, n_102);
  nand g364 (n_452, n_103, n_102);
  nand g365 (n_453, n_101, n_103);
  nand g366 (out_0[6], n_451, n_452, n_453);
  xor g367 (n_118, n_104, n_105);
  and g368 (n_152, n_104, n_105);
  xor g369 (n_454, n_106, n_107);
  xor g370 (n_123, n_454, n_108);
  nand g371 (n_455, n_106, n_107);
  nand g372 (n_456, n_108, n_107);
  nand g373 (n_457, n_106, n_108);
  nand g374 (n_154, n_455, n_456, n_457);
  xor g375 (n_458, n_109, n_110);
  xor g376 (n_125, n_458, n_111);
  nand g377 (n_459, n_109, n_110);
  nand g378 (n_460, n_111, n_110);
  nand g379 (n_461, n_109, n_111);
  nand g380 (n_157, n_459, n_460, n_461);
  xor g381 (n_462, n_112, n_113);
  xor g382 (n_126, n_462, n_114);
  nand g383 (n_463, n_112, n_113);
  nand g384 (n_464, n_114, n_113);
  nand g385 (n_465, n_112, n_114);
  nand g386 (n_155, n_463, n_464, n_465);
  xor g387 (n_466, n_115, n_116);
  xor g388 (n_124, n_466, n_117);
  nand g389 (n_467, n_115, n_116);
  nand g390 (n_468, n_117, n_116);
  nand g391 (n_469, n_115, n_117);
  nand g392 (n_156, n_467, n_468, n_469);
  xor g393 (n_470, n_118, n_119);
  xor g394 (n_128, n_470, n_120);
  nand g395 (n_471, n_118, n_119);
  nand g396 (n_472, n_120, n_119);
  nand g397 (n_473, n_118, n_120);
  nand g398 (n_163, n_471, n_472, n_473);
  xor g399 (n_474, n_121, n_122);
  xor g400 (n_129, n_474, n_123);
  nand g401 (n_475, n_121, n_122);
  nand g402 (n_476, n_123, n_122);
  nand g403 (n_477, n_121, n_123);
  nand g404 (n_165, n_475, n_476, n_477);
  xor g405 (n_478, n_124, n_125);
  xor g406 (n_131, n_478, n_126);
  nand g407 (n_479, n_124, n_125);
  nand g408 (n_480, n_126, n_125);
  nand g409 (n_481, n_124, n_126);
  nand g410 (n_164, n_479, n_480, n_481);
  xor g411 (n_482, n_127, n_128);
  xor g412 (n_133, n_482, n_129);
  nand g413 (n_483, n_127, n_128);
  nand g414 (n_484, n_129, n_128);
  nand g415 (n_485, n_127, n_129);
  nand g416 (n_169, n_483, n_484, n_485);
  xor g417 (n_486, n_130, n_131);
  xor g418 (n_135, n_486, n_132);
  nand g419 (n_487, n_130, n_131);
  nand g420 (n_488, n_132, n_131);
  nand g421 (n_489, n_130, n_132);
  nand g422 (n_172, n_487, n_488, n_489);
  xor g423 (n_490, n_133, n_134);
  xor g424 (out_1[6], n_490, n_135);
  nand g425 (n_491, n_133, n_134);
  nand g426 (n_492, n_135, n_134);
  nand g427 (n_493, n_133, n_135);
  nand g428 (out_0[7], n_491, n_492, n_493);
  xor g429 (n_153, n_136, n_137);
  and g430 (n_189, n_136, n_137);
  xor g431 (n_494, n_138, n_139);
  xor g432 (n_159, n_494, n_140);
  nand g433 (n_495, n_138, n_139);
  nand g434 (n_496, n_140, n_139);
  nand g435 (n_497, n_138, n_140);
  nand g436 (n_190, n_495, n_496, n_497);
  xor g437 (n_498, n_141, n_142);
  xor g438 (n_160, n_498, n_143);
  nand g439 (n_499, n_141, n_142);
  nand g440 (n_500, n_143, n_142);
  nand g441 (n_501, n_141, n_143);
  nand g442 (n_191, n_499, n_500, n_501);
  xor g443 (n_502, n_144, n_145);
  xor g444 (n_158, n_502, n_146);
  nand g445 (n_503, n_144, n_145);
  nand g446 (n_504, n_146, n_145);
  nand g447 (n_505, n_144, n_146);
  nand g448 (n_192, n_503, n_504, n_505);
  xor g449 (n_506, n_147, n_148);
  xor g450 (n_161, n_506, n_149);
  nand g451 (n_507, n_147, n_148);
  nand g452 (n_508, n_149, n_148);
  nand g453 (n_509, n_147, n_149);
  nand g454 (n_193, n_507, n_508, n_509);
  xor g455 (n_510, n_150, n_151);
  xor g456 (n_162, n_510, n_152);
  nand g457 (n_511, n_150, n_151);
  nand g458 (n_512, n_152, n_151);
  nand g459 (n_513, n_150, n_152);
  nand g460 (n_198, n_511, n_512, n_513);
  xor g461 (n_514, n_153, n_154);
  xor g462 (n_166, n_514, n_155);
  nand g463 (n_515, n_153, n_154);
  nand g464 (n_516, n_155, n_154);
  nand g465 (n_517, n_153, n_155);
  nand g466 (n_200, n_515, n_516, n_517);
  xor g467 (n_518, n_156, n_157);
  xor g468 (n_167, n_518, n_158);
  nand g469 (n_519, n_156, n_157);
  nand g470 (n_520, n_158, n_157);
  nand g471 (n_521, n_156, n_158);
  nand g472 (n_201, n_519, n_520, n_521);
  xor g473 (n_522, n_159, n_160);
  xor g474 (n_168, n_522, n_161);
  nand g475 (n_523, n_159, n_160);
  nand g476 (n_524, n_161, n_160);
  nand g477 (n_525, n_159, n_161);
  nand g478 (n_202, n_523, n_524, n_525);
  xor g479 (n_526, n_162, n_163);
  xor g480 (n_170, n_526, n_164);
  nand g481 (n_527, n_162, n_163);
  nand g482 (n_528, n_164, n_163);
  nand g483 (n_529, n_162, n_164);
  nand g484 (n_207, n_527, n_528, n_529);
  xor g485 (n_530, n_165, n_166);
  xor g486 (n_171, n_530, n_167);
  nand g487 (n_531, n_165, n_166);
  nand g488 (n_532, n_167, n_166);
  nand g489 (n_533, n_165, n_167);
  nand g490 (n_206, n_531, n_532, n_533);
  xor g491 (n_534, n_168, n_169);
  xor g492 (n_173, n_534, n_170);
  nand g493 (n_535, n_168, n_169);
  nand g494 (n_536, n_170, n_169);
  nand g495 (n_537, n_168, n_170);
  nand g496 (n_210, n_535, n_536, n_537);
  xor g497 (n_538, n_171, n_172);
  xor g498 (out_1[7], n_538, n_173);
  nand g499 (n_539, n_171, n_172);
  nand g500 (n_540, n_173, n_172);
  nand g501 (n_541, n_171, n_173);
  nand g502 (out_0[8], n_539, n_540, n_541);
  xor g503 (n_188, n_174, n_175);
  and g504 (n_225, n_174, n_175);
  xor g505 (n_542, n_176, n_177);
  xor g506 (n_194, n_542, n_178);
  nand g507 (n_543, n_176, n_177);
  nand g508 (n_544, n_178, n_177);
  nand g509 (n_545, n_176, n_178);
  nand g510 (n_228, n_543, n_544, n_545);
  xor g511 (n_546, n_179, n_180);
  xor g512 (n_196, n_546, n_181);
  nand g513 (n_547, n_179, n_180);
  nand g514 (n_548, n_181, n_180);
  nand g515 (n_549, n_179, n_181);
  nand g516 (n_229, n_547, n_548, n_549);
  xor g517 (n_550, n_182, n_183);
  xor g518 (n_195, n_550, n_184);
  nand g519 (n_551, n_182, n_183);
  nand g520 (n_552, n_184, n_183);
  nand g521 (n_553, n_182, n_184);
  nand g522 (n_226, n_551, n_552, n_553);
  xor g523 (n_554, n_185, n_186);
  xor g524 (n_197, n_554, n_187);
  nand g525 (n_555, n_185, n_186);
  nand g526 (n_556, n_187, n_186);
  nand g527 (n_557, n_185, n_187);
  nand g528 (n_227, n_555, n_556, n_557);
  xor g529 (n_558, n_188, n_189);
  xor g530 (n_199, n_558, n_190);
  nand g531 (n_559, n_188, n_189);
  nand g532 (n_560, n_190, n_189);
  nand g533 (n_561, n_188, n_190);
  nand g534 (n_234, n_559, n_560, n_561);
  xor g535 (n_562, n_191, n_192);
  xor g536 (n_203, n_562, n_193);
  nand g537 (n_563, n_191, n_192);
  nand g538 (n_564, n_193, n_192);
  nand g539 (n_565, n_191, n_193);
  nand g540 (n_235, n_563, n_564, n_565);
  xor g541 (n_566, n_194, n_195);
  xor g542 (n_204, n_566, n_196);
  nand g543 (n_567, n_194, n_195);
  nand g544 (n_568, n_196, n_195);
  nand g545 (n_569, n_194, n_196);
  nand g546 (n_236, n_567, n_568, n_569);
  xor g547 (n_570, n_197, n_198);
  xor g548 (n_205, n_570, n_199);
  nand g549 (n_571, n_197, n_198);
  nand g550 (n_572, n_199, n_198);
  nand g551 (n_573, n_197, n_199);
  nand g552 (n_239, n_571, n_572, n_573);
  xor g553 (n_574, n_200, n_201);
  xor g554 (n_208, n_574, n_202);
  nand g555 (n_575, n_200, n_201);
  nand g556 (n_576, n_202, n_201);
  nand g557 (n_577, n_200, n_202);
  nand g558 (n_240, n_575, n_576, n_577);
  xor g559 (n_578, n_203, n_204);
  xor g560 (n_209, n_578, n_205);
  nand g561 (n_579, n_203, n_204);
  nand g562 (n_580, n_205, n_204);
  nand g563 (n_581, n_203, n_205);
  nand g564 (n_243, n_579, n_580, n_581);
  xor g565 (n_582, n_206, n_207);
  xor g566 (n_211, n_582, n_208);
  nand g567 (n_583, n_206, n_207);
  nand g568 (n_584, n_208, n_207);
  nand g569 (n_585, n_206, n_208);
  nand g570 (n_245, n_583, n_584, n_585);
  xor g571 (n_586, n_209, n_210);
  xor g572 (out_1[8], n_586, n_211);
  nand g573 (n_587, n_209, n_210);
  nand g574 (n_588, n_211, n_210);
  nand g575 (n_589, n_209, n_211);
  nand g576 (out_0[9], n_587, n_588, n_589);
  xor g577 (n_224, n_212, n_213);
  and g578 (n_257, n_212, n_213);
  xor g579 (n_590, n_214, n_215);
  xor g580 (n_231, n_590, n_216);
  nand g581 (n_591, n_214, n_215);
  nand g582 (n_592, n_216, n_215);
  nand g583 (n_593, n_214, n_216);
  nand g584 (n_258, n_591, n_592, n_593);
  xor g585 (n_594, n_217, n_218);
  xor g586 (n_232, n_594, n_219);
  nand g587 (n_595, n_217, n_218);
  nand g588 (n_596, n_219, n_218);
  nand g589 (n_597, n_217, n_219);
  nand g590 (n_259, n_595, n_596, n_597);
  xor g591 (n_598, n_220, n_221);
  xor g592 (n_230, n_598, n_222);
  nand g593 (n_599, n_220, n_221);
  nand g594 (n_600, n_222, n_221);
  nand g595 (n_601, n_220, n_222);
  nand g596 (n_260, n_599, n_600, n_601);
  xor g597 (n_602, n_223, n_224);
  xor g598 (n_233, n_602, n_225);
  nand g599 (n_603, n_223, n_224);
  nand g600 (n_604, n_225, n_224);
  nand g601 (n_605, n_223, n_225);
  nand g602 (n_264, n_603, n_604, n_605);
  xor g603 (n_606, n_226, n_227);
  xor g604 (n_237, n_606, n_228);
  nand g605 (n_607, n_226, n_227);
  nand g606 (n_608, n_228, n_227);
  nand g607 (n_609, n_226, n_228);
  nand g608 (n_265, n_607, n_608, n_609);
  xor g609 (n_610, n_229, n_230);
  xor g610 (n_238, n_610, n_231);
  nand g611 (n_611, n_229, n_230);
  nand g612 (n_612, n_231, n_230);
  nand g613 (n_613, n_229, n_231);
  nand g614 (n_267, n_611, n_612, n_613);
  xor g615 (n_614, n_232, n_233);
  xor g616 (n_241, n_614, n_234);
  nand g617 (n_615, n_232, n_233);
  nand g618 (n_616, n_234, n_233);
  nand g619 (n_617, n_232, n_234);
  nand g620 (n_270, n_615, n_616, n_617);
  xor g621 (n_618, n_235, n_236);
  xor g622 (n_242, n_618, n_237);
  nand g623 (n_619, n_235, n_236);
  nand g624 (n_620, n_237, n_236);
  nand g625 (n_621, n_235, n_237);
  nand g626 (n_272, n_619, n_620, n_621);
  xor g627 (n_622, n_238, n_239);
  xor g628 (n_244, n_622, n_240);
  nand g629 (n_623, n_238, n_239);
  nand g630 (n_624, n_240, n_239);
  nand g631 (n_625, n_238, n_240);
  nand g632 (n_274, n_623, n_624, n_625);
  xor g633 (n_626, n_241, n_242);
  xor g634 (n_246, n_626, n_243);
  nand g635 (n_627, n_241, n_242);
  nand g636 (n_628, n_243, n_242);
  nand g637 (n_629, n_241, n_243);
  nand g638 (n_276, n_627, n_628, n_629);
  xor g639 (n_630, n_244, n_245);
  xor g640 (out_1[9], n_630, n_246);
  nand g641 (n_631, n_244, n_245);
  nand g642 (n_632, n_246, n_245);
  nand g643 (n_633, n_244, n_246);
  nand g644 (out_0[10], n_631, n_632, n_633);
  xor g645 (n_634, n_247, n_248);
  xor g646 (n_263, n_634, n_249);
  nand g647 (n_635, n_247, n_248);
  nand g648 (n_636, n_249, n_248);
  nand g649 (n_637, n_247, n_249);
  nand g650 (n_285, n_635, n_636, n_637);
  xor g651 (n_638, n_250, n_251);
  xor g652 (n_261, n_638, n_252);
  nand g653 (n_639, n_250, n_251);
  nand g654 (n_640, n_252, n_251);
  nand g655 (n_641, n_250, n_252);
  nand g656 (n_286, n_639, n_640, n_641);
  xor g657 (n_642, n_253, n_254);
  xor g658 (n_262, n_642, n_255);
  nand g659 (n_643, n_253, n_254);
  nand g660 (n_644, n_255, n_254);
  nand g661 (n_645, n_253, n_255);
  nand g662 (n_287, n_643, n_644, n_645);
  xor g663 (n_646, n_256, n_257);
  xor g664 (n_266, n_646, n_258);
  nand g665 (n_647, n_256, n_257);
  nand g666 (n_648, n_258, n_257);
  nand g667 (n_649, n_256, n_258);
  nand g668 (n_291, n_647, n_648, n_649);
  xor g669 (n_650, n_259, n_260);
  xor g670 (n_268, n_650, n_261);
  nand g671 (n_651, n_259, n_260);
  nand g672 (n_652, n_261, n_260);
  nand g673 (n_653, n_259, n_261);
  nand g674 (n_293, n_651, n_652, n_653);
  xor g675 (n_654, n_262, n_263);
  xor g676 (n_269, n_654, n_264);
  nand g677 (n_655, n_262, n_263);
  nand g678 (n_656, n_264, n_263);
  nand g679 (n_657, n_262, n_264);
  nand g680 (n_294, n_655, n_656, n_657);
  xor g681 (n_658, n_265, n_266);
  xor g682 (n_271, n_658, n_267);
  nand g683 (n_659, n_265, n_266);
  nand g684 (n_660, n_267, n_266);
  nand g685 (n_661, n_265, n_267);
  nand g686 (n_296, n_659, n_660, n_661);
  xor g687 (n_662, n_268, n_269);
  xor g688 (n_273, n_662, n_270);
  nand g689 (n_663, n_268, n_269);
  nand g690 (n_664, n_270, n_269);
  nand g691 (n_665, n_268, n_270);
  nand g692 (n_298, n_663, n_664, n_665);
  xor g693 (n_666, n_271, n_272);
  xor g694 (n_275, n_666, n_273);
  nand g695 (n_667, n_271, n_272);
  nand g696 (n_668, n_273, n_272);
  nand g697 (n_669, n_271, n_273);
  nand g698 (n_300, n_667, n_668, n_669);
  xor g699 (n_670, n_274, n_275);
  xor g700 (out_1[10], n_670, n_276);
  nand g701 (n_671, n_274, n_275);
  nand g702 (n_672, n_276, n_275);
  nand g703 (n_673, n_274, n_276);
  nand g704 (out_0[11], n_671, n_672, n_673);
  xor g705 (n_674, n_277, n_278);
  xor g706 (n_288, n_674, n_279);
  nand g707 (n_675, n_277, n_278);
  nand g708 (n_676, n_279, n_278);
  nand g709 (n_677, n_277, n_279);
  nand g710 (n_308, n_675, n_676, n_677);
  xor g711 (n_678, n_280, n_281);
  xor g712 (n_289, n_678, n_282);
  nand g713 (n_679, n_280, n_281);
  nand g714 (n_680, n_282, n_281);
  nand g715 (n_681, n_280, n_282);
  nand g716 (n_307, n_679, n_680, n_681);
  xor g717 (n_682, n_283, n_284);
  xor g718 (n_290, n_682, n_285);
  nand g719 (n_683, n_283, n_284);
  nand g720 (n_684, n_285, n_284);
  nand g721 (n_685, n_283, n_285);
  nand g722 (n_311, n_683, n_684, n_685);
  xor g723 (n_686, n_286, n_287);
  xor g724 (n_292, n_686, n_288);
  nand g725 (n_687, n_286, n_287);
  nand g726 (n_688, n_288, n_287);
  nand g727 (n_689, n_286, n_288);
  nand g728 (n_313, n_687, n_688, n_689);
  xor g729 (n_690, n_289, n_290);
  xor g730 (n_295, n_690, n_291);
  nand g731 (n_691, n_289, n_290);
  nand g732 (n_692, n_291, n_290);
  nand g733 (n_693, n_289, n_291);
  nand g734 (n_314, n_691, n_692, n_693);
  xor g735 (n_694, n_292, n_293);
  xor g736 (n_297, n_694, n_294);
  nand g737 (n_695, n_292, n_293);
  nand g738 (n_696, n_294, n_293);
  nand g739 (n_697, n_292, n_294);
  nand g740 (n_316, n_695, n_696, n_697);
  xor g741 (n_698, n_295, n_296);
  xor g742 (n_299, n_698, n_297);
  nand g743 (n_699, n_295, n_296);
  nand g744 (n_700, n_297, n_296);
  nand g745 (n_701, n_295, n_297);
  nand g746 (n_318, n_699, n_700, n_701);
  xor g747 (n_702, n_298, n_299);
  xor g748 (out_1[11], n_702, n_300);
  nand g749 (n_703, n_298, n_299);
  nand g750 (n_704, n_300, n_299);
  nand g751 (n_705, n_298, n_300);
  nand g752 (out_1[12], n_703, n_704, n_705);
  xor g753 (n_706, n_301, n_302);
  xor g754 (n_310, n_706, n_303);
  nand g755 (n_707, n_301, n_302);
  nand g756 (n_708, n_303, n_302);
  nand g757 (n_709, n_301, n_303);
  nand g758 (n_323, n_707, n_708, n_709);
  xor g759 (n_710, n_304, n_305);
  xor g760 (n_309, n_710, n_306);
  nand g761 (n_711, n_304, n_305);
  nand g762 (n_712, n_306, n_305);
  nand g763 (n_713, n_304, n_306);
  nand g764 (n_324, n_711, n_712, n_713);
  xor g765 (n_714, n_307, n_308);
  xor g766 (n_312, n_714, n_309);
  nand g767 (n_715, n_307, n_308);
  nand g768 (n_716, n_309, n_308);
  nand g769 (n_717, n_307, n_309);
  nand g770 (n_327, n_715, n_716, n_717);
  xor g771 (n_718, n_310, n_311);
  xor g772 (n_315, n_718, n_312);
  nand g773 (n_719, n_310, n_311);
  nand g774 (n_720, n_312, n_311);
  nand g775 (n_721, n_310, n_312);
  nand g776 (n_328, n_719, n_720, n_721);
  xor g777 (n_722, n_313, n_314);
  xor g778 (n_317, n_722, n_315);
  nand g779 (n_723, n_313, n_314);
  nand g780 (n_724, n_315, n_314);
  nand g781 (n_725, n_313, n_315);
  nand g782 (n_330, n_723, n_724, n_725);
  xor g783 (n_726, n_316, n_317);
  xor g784 (out_0[12], n_726, n_318);
  nand g785 (n_727, n_316, n_317);
  nand g786 (n_728, n_318, n_317);
  nand g787 (n_729, n_316, n_318);
  nand g788 (out_1[13], n_727, n_728, n_729);
  xor g789 (n_730, n_319, n_320);
  xor g790 (n_325, n_730, n_321);
  nand g791 (n_731, n_319, n_320);
  nand g792 (n_732, n_321, n_320);
  nand g793 (n_733, n_319, n_321);
  nand g794 (n_333, n_731, n_732, n_733);
  xor g795 (n_734, n_322, n_323);
  xor g796 (n_326, n_734, n_324);
  nand g797 (n_735, n_322, n_323);
  nand g798 (n_736, n_324, n_323);
  nand g799 (n_737, n_322, n_324);
  nand g800 (n_334, n_735, n_736, n_737);
  xor g801 (n_738, n_325, n_326);
  xor g802 (n_329, n_738, n_327);
  nand g803 (n_739, n_325, n_326);
  nand g804 (n_740, n_327, n_326);
  nand g805 (n_741, n_325, n_327);
  nand g806 (n_336, n_739, n_740, n_741);
  xor g807 (n_742, n_328, n_329);
  xor g808 (out_0[13], n_742, n_330);
  nand g809 (n_743, n_328, n_329);
  nand g810 (n_744, n_330, n_329);
  nand g811 (n_745, n_328, n_330);
  nand g812 (out_1[14], n_743, n_744, n_745);
  xor g813 (n_746, n_331, n_332);
  xor g814 (n_335, n_746, n_333);
  nand g815 (n_747, n_331, n_332);
  nand g816 (n_748, n_333, n_332);
  nand g817 (n_749, n_331, n_333);
  nand g818 (out_0[15], n_747, n_748, n_749);
  xor g819 (n_750, n_334, n_335);
  xor g820 (out_0[14], n_750, n_336);
  nand g821 (n_751, n_334, n_335);
  nand g822 (n_752, n_336, n_335);
  nand g823 (n_753, n_334, n_336);
  nand g824 (out_1[15], n_751, n_752, n_753);
endmodule

module csa_tree_GENERIC(in_0, in_1, in_2, in_3, out_0, out_1);
  input [7:0] in_0, in_1, in_2, in_3;
  output [16:0] out_0, out_1;
  wire [7:0] in_0, in_1, in_2, in_3;
  wire [16:0] out_0, out_1;
  csa_tree_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2 (in_2),
       .in_3 (in_3), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_271_GENERIC_REAL(in_0, in_1, in_2, in_3, out_0, out_1,
     out_2);
// synthesis_equation "assign out_0 = ( ( in_2 + in_3 ) + ( in_0 * in_1 )  )  ; assign out_1 = 17'b0; assign out_2 = 1'b0;"
  input [16:0] in_0, in_2, in_3;
  input [7:0] in_1;
  output [16:0] out_0, out_1;
  output out_2;
  wire [16:0] in_0, in_2, in_3;
  wire [7:0] in_1;
  wire [16:0] out_0, out_1;
  wire out_2;
  wire n_27, n_30, n_32, n_33, n_34, n_35, n_37, n_39;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_74, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_86, n_87, n_88, n_89, n_90, n_91, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_135, n_136, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251;
  wire n_252, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602;
  wire n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610;
  wire n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618;
  wire n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642;
  wire n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650;
  wire n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682;
  wire n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698;
  wire n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706;
  wire n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714;
  wire n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_725;
  wire n_729, n_733, n_737, n_741, n_745;
  assign out_2 = in_2[0];
  assign out_0[0] = in_3[0];
  and g1 (out_1[0], in_0[0], in_1[0]);
  and g2 (out_0[1], in_0[1], in_1[0]);
  and g3 (out_0[2], in_0[2], in_1[0]);
  and g4 (n_42, in_0[3], in_1[0]);
  and g5 (n_55, in_0[4], in_1[0]);
  and g6 (n_69, in_0[5], in_1[0]);
  and g7 (n_85, in_0[6], in_1[0]);
  and g8 (n_106, in_0[7], in_1[0]);
  and g9 (n_128, in_0[8], in_1[0]);
  and g10 (n_150, in_0[9], in_1[0]);
  and g11 (n_173, in_0[10], in_1[0]);
  and g12 (n_196, in_0[11], in_1[0]);
  and g13 (n_220, in_0[12], in_1[0]);
  and g14 (n_245, in_0[13], in_1[0]);
  and g15 (n_266, in_0[14], in_1[0]);
  and g16 (n_289, in_0[15], in_1[0]);
  and g17 (n_314, in_0[16], in_1[0]);
  and g18 (n_27, in_0[0], in_1[1]);
  and g19 (n_32, in_0[1], in_1[1]);
  and g20 (n_41, in_0[2], in_1[1]);
  and g21 (n_51, in_0[3], in_1[1]);
  and g22 (n_66, in_0[4], in_1[1]);
  and g23 (n_84, in_0[5], in_1[1]);
  and g24 (n_103, in_0[6], in_1[1]);
  and g25 (n_125, in_0[7], in_1[1]);
  and g26 (n_149, in_0[8], in_1[1]);
  and g27 (n_172, in_0[9], in_1[1]);
  and g28 (n_194, in_0[10], in_1[1]);
  and g29 (n_219, in_0[11], in_1[1]);
  and g30 (n_242, in_0[12], in_1[1]);
  and g31 (n_267, in_0[13], in_1[1]);
  and g32 (n_287, in_0[14], in_1[1]);
  and g33 (n_310, in_0[15], in_1[1]);
  and g34 (n_30, in_0[0], in_1[2]);
  and g35 (n_37, in_0[1], in_1[2]);
  and g36 (n_49, in_0[2], in_1[2]);
  and g37 (n_63, in_0[3], in_1[2]);
  and g38 (n_80, in_0[4], in_1[2]);
  and g39 (n_101, in_0[5], in_1[2]);
  and g40 (n_121, in_0[6], in_1[2]);
  and g41 (n_147, in_0[7], in_1[2]);
  and g42 (n_170, in_0[8], in_1[2]);
  and g43 (n_193, in_0[9], in_1[2]);
  and g44 (n_215, in_0[10], in_1[2]);
  and g45 (n_239, in_0[11], in_1[2]);
  and g46 (n_263, in_0[12], in_1[2]);
  and g47 (n_288, in_0[13], in_1[2]);
  and g48 (n_306, in_0[14], in_1[2]);
  and g49 (n_35, in_0[0], in_1[3]);
  and g50 (n_45, in_0[1], in_1[3]);
  and g51 (n_61, in_0[2], in_1[3]);
  and g52 (n_77, in_0[3], in_1[3]);
  and g53 (n_98, in_0[4], in_1[3]);
  and g54 (n_120, in_0[5], in_1[3]);
  and g55 (n_143, in_0[6], in_1[3]);
  and g56 (n_167, in_0[7], in_1[3]);
  and g57 (n_191, in_0[8], in_1[3]);
  and g58 (n_214, in_0[9], in_1[3]);
  and g59 (n_238, in_0[10], in_1[3]);
  and g60 (n_262, in_0[11], in_1[3]);
  and g61 (n_286, in_0[12], in_1[3]);
  and g62 (n_307, in_0[13], in_1[3]);
  and g63 (n_44, in_0[0], in_1[4]);
  and g64 (n_57, in_0[1], in_1[4]);
  and g65 (n_74, in_0[2], in_1[4]);
  and g66 (n_94, in_0[3], in_1[4]);
  and g67 (n_118, in_0[4], in_1[4]);
  and g68 (n_141, in_0[5], in_1[4]);
  and g69 (n_165, in_0[6], in_1[4]);
  and g70 (n_189, in_0[7], in_1[4]);
  and g71 (n_213, in_0[8], in_1[4]);
  and g72 (n_236, in_0[9], in_1[4]);
  and g73 (n_260, in_0[10], in_1[4]);
  and g74 (n_284, in_0[11], in_1[4]);
  and g75 (n_305, in_0[12], in_1[4]);
  and g76 (n_56, in_0[0], in_1[5]);
  and g77 (n_72, in_0[1], in_1[5]);
  and g78 (n_91, in_0[2], in_1[5]);
  and g79 (n_112, in_0[3], in_1[5]);
  and g80 (n_138, in_0[4], in_1[5]);
  and g81 (n_163, in_0[5], in_1[5]);
  and g82 (n_187, in_0[6], in_1[5]);
  and g83 (n_211, in_0[7], in_1[5]);
  and g84 (n_235, in_0[8], in_1[5]);
  and g85 (n_258, in_0[9], in_1[5]);
  and g86 (n_281, in_0[10], in_1[5]);
  and g87 (n_304, in_0[11], in_1[5]);
  and g88 (n_71, in_0[0], in_1[6]);
  and g89 (n_90, in_0[1], in_1[6]);
  and g90 (n_111, in_0[2], in_1[6]);
  and g91 (n_135, in_0[3], in_1[6]);
  and g92 (n_160, in_0[4], in_1[6]);
  and g93 (n_184, in_0[5], in_1[6]);
  and g94 (n_208, in_0[6], in_1[6]);
  and g95 (n_232, in_0[7], in_1[6]);
  and g96 (n_256, in_0[8], in_1[6]);
  and g97 (n_280, in_0[9], in_1[6]);
  and g98 (n_302, in_0[10], in_1[6]);
  and g99 (n_89, in_0[0], in_1[7]);
  and g100 (n_110, in_0[1], in_1[7]);
  and g101 (n_133, in_0[2], in_1[7]);
  and g102 (n_157, in_0[3], in_1[7]);
  and g103 (n_183, in_0[4], in_1[7]);
  and g104 (n_207, in_0[5], in_1[7]);
  and g105 (n_231, in_0[6], in_1[7]);
  and g106 (n_255, in_0[7], in_1[7]);
  and g107 (n_279, in_0[8], in_1[7]);
  and g108 (n_301, in_0[9], in_1[7]);
  xor g208 (n_357, in_2[1], n_27);
  xor g209 (out_1[1], n_357, in_3[1]);
  nand g210 (n_358, in_2[1], n_27);
  nand g211 (n_359, in_3[1], n_27);
  nand g212 (n_360, in_2[1], in_3[1]);
  nand g213 (n_33, n_358, n_359, n_360);
  xor g214 (n_361, in_2[2], n_30);
  xor g215 (n_34, n_361, in_3[2]);
  nand g216 (n_362, in_2[2], n_30);
  nand g217 (n_363, in_3[2], n_30);
  nand g218 (n_364, in_2[2], in_3[2]);
  nand g219 (n_39, n_362, n_363, n_364);
  xor g220 (n_365, n_32, n_33);
  xor g221 (out_1[2], n_365, n_34);
  nand g222 (n_366, n_32, n_33);
  nand g223 (n_367, n_34, n_33);
  nand g224 (n_368, n_32, n_34);
  nand g225 (n_43, n_366, n_367, n_368);
  xor g226 (n_369, n_35, in_2[3]);
  xor g227 (n_40, n_369, n_37);
  nand g228 (n_370, n_35, in_2[3]);
  nand g229 (n_371, n_37, in_2[3]);
  nand g230 (n_372, n_35, n_37);
  nand g231 (n_48, n_370, n_371, n_372);
  xor g232 (n_373, in_3[3], n_39);
  xor g233 (out_0[3], n_373, n_40);
  nand g234 (n_374, in_3[3], n_39);
  nand g235 (n_375, n_40, n_39);
  nand g236 (n_376, in_3[3], n_40);
  nand g237 (n_52, n_374, n_375, n_376);
  xor g238 (n_377, n_41, n_42);
  xor g239 (out_1[3], n_377, n_43);
  nand g240 (n_378, n_41, n_42);
  nand g241 (n_379, n_43, n_42);
  nand g242 (n_380, n_41, n_43);
  nand g243 (n_54, n_378, n_379, n_380);
  xor g244 (n_381, n_44, n_45);
  xor g245 (n_50, n_381, in_2[4]);
  nand g246 (n_382, n_44, n_45);
  nand g247 (n_383, in_2[4], n_45);
  nand g248 (n_384, n_44, in_2[4]);
  nand g249 (n_60, n_382, n_383, n_384);
  xor g250 (n_385, in_3[4], n_48);
  xor g251 (n_53, n_385, n_49);
  nand g252 (n_386, in_3[4], n_48);
  nand g253 (n_387, n_49, n_48);
  nand g254 (n_388, in_3[4], n_49);
  nand g255 (n_64, n_386, n_387, n_388);
  xor g256 (n_389, n_50, n_51);
  xor g257 (out_0[4], n_389, n_52);
  nand g258 (n_390, n_50, n_51);
  nand g259 (n_391, n_52, n_51);
  nand g260 (n_392, n_50, n_52);
  nand g261 (n_67, n_390, n_391, n_392);
  xor g262 (n_393, n_53, n_54);
  xor g263 (out_1[4], n_393, n_55);
  nand g264 (n_394, n_53, n_54);
  nand g265 (n_395, n_55, n_54);
  nand g266 (n_396, n_53, n_55);
  nand g267 (n_70, n_394, n_395, n_396);
  xor g268 (n_397, n_56, n_57);
  xor g269 (n_62, n_397, in_2[5]);
  nand g270 (n_398, n_56, n_57);
  nand g271 (n_399, in_2[5], n_57);
  nand g272 (n_400, n_56, in_2[5]);
  nand g273 (n_76, n_398, n_399, n_400);
  xor g274 (n_401, in_3[5], n_60);
  xor g275 (n_65, n_401, n_61);
  nand g276 (n_402, in_3[5], n_60);
  nand g277 (n_403, n_61, n_60);
  nand g278 (n_404, in_3[5], n_61);
  nand g279 (n_78, n_402, n_403, n_404);
  xor g280 (n_405, n_62, n_63);
  xor g281 (n_68, n_405, n_64);
  nand g282 (n_406, n_62, n_63);
  nand g283 (n_407, n_64, n_63);
  nand g284 (n_408, n_62, n_64);
  nand g285 (n_82, n_406, n_407, n_408);
  xor g286 (n_409, n_65, n_66);
  xor g287 (out_0[5], n_409, n_67);
  nand g288 (n_410, n_65, n_66);
  nand g289 (n_411, n_67, n_66);
  nand g290 (n_412, n_65, n_67);
  nand g291 (n_86, n_410, n_411, n_412);
  xor g292 (n_413, n_68, n_69);
  xor g293 (out_1[5], n_413, n_70);
  nand g294 (n_414, n_68, n_69);
  nand g295 (n_415, n_70, n_69);
  nand g296 (n_416, n_68, n_70);
  nand g297 (out_0[6], n_414, n_415, n_416);
  xor g298 (n_417, n_71, n_72);
  xor g299 (n_79, n_417, in_2[6]);
  nand g300 (n_418, n_71, n_72);
  nand g301 (n_419, in_2[6], n_72);
  nand g302 (n_420, n_71, in_2[6]);
  nand g303 (n_96, n_418, n_419, n_420);
  xor g304 (n_421, n_74, in_3[6]);
  xor g305 (n_81, n_421, n_76);
  nand g306 (n_422, n_74, in_3[6]);
  nand g307 (n_423, n_76, in_3[6]);
  nand g308 (n_424, n_74, n_76);
  nand g309 (n_97, n_422, n_423, n_424);
  xor g310 (n_425, n_77, n_78);
  xor g311 (n_83, n_425, n_79);
  nand g312 (n_426, n_77, n_78);
  nand g313 (n_427, n_79, n_78);
  nand g314 (n_428, n_77, n_79);
  nand g315 (n_99, n_426, n_427, n_428);
  xor g316 (n_429, n_80, n_81);
  xor g317 (n_87, n_429, n_82);
  nand g318 (n_430, n_80, n_81);
  nand g319 (n_431, n_82, n_81);
  nand g320 (n_432, n_80, n_82);
  nand g321 (n_104, n_430, n_431, n_432);
  xor g322 (n_433, n_83, n_84);
  xor g323 (n_88, n_433, n_85);
  nand g324 (n_434, n_83, n_84);
  nand g325 (n_435, n_85, n_84);
  nand g326 (n_436, n_83, n_85);
  nand g327 (n_107, n_434, n_435, n_436);
  xor g328 (n_437, n_86, n_87);
  xor g329 (out_1[6], n_437, n_88);
  nand g330 (n_438, n_86, n_87);
  nand g331 (n_439, n_88, n_87);
  nand g332 (n_440, n_86, n_88);
  nand g333 (n_109, n_438, n_439, n_440);
  xor g334 (n_441, n_89, n_90);
  xor g335 (n_95, n_441, n_91);
  nand g336 (n_442, n_89, n_90);
  nand g337 (n_443, n_91, n_90);
  nand g338 (n_444, n_89, n_91);
  nand g339 (n_116, n_442, n_443, n_444);
  xor g340 (n_445, in_2[7], in_3[7]);
  xor g341 (n_100, n_445, n_94);
  nand g342 (n_446, in_2[7], in_3[7]);
  nand g343 (n_447, n_94, in_3[7]);
  nand g344 (n_448, in_2[7], n_94);
  nand g345 (n_117, n_446, n_447, n_448);
  xor g346 (n_449, n_95, n_96);
  xor g347 (n_102, n_449, n_97);
  nand g348 (n_450, n_95, n_96);
  nand g349 (n_451, n_97, n_96);
  nand g350 (n_452, n_95, n_97);
  nand g351 (n_122, n_450, n_451, n_452);
  xor g352 (n_453, n_98, n_99);
  xor g353 (n_105, n_453, n_100);
  nand g354 (n_454, n_98, n_99);
  nand g355 (n_455, n_100, n_99);
  nand g356 (n_456, n_98, n_100);
  nand g357 (n_124, n_454, n_455, n_456);
  xor g358 (n_457, n_101, n_102);
  xor g359 (n_108, n_457, n_103);
  nand g360 (n_458, n_101, n_102);
  nand g361 (n_459, n_103, n_102);
  nand g362 (n_460, n_101, n_103);
  nand g363 (n_127, n_458, n_459, n_460);
  xor g364 (n_461, n_104, n_105);
  xor g365 (out_0[7], n_461, n_106);
  nand g366 (n_462, n_104, n_105);
  nand g367 (n_463, n_106, n_105);
  nand g368 (n_464, n_104, n_106);
  nand g369 (n_130, n_462, n_463, n_464);
  xor g370 (n_465, n_107, n_108);
  xor g371 (out_1[7], n_465, n_109);
  nand g372 (n_466, n_107, n_108);
  nand g373 (n_467, n_109, n_108);
  nand g374 (n_468, n_107, n_109);
  nand g375 (out_0[8], n_466, n_467, n_468);
  xor g376 (n_113, n_110, n_111);
  and g377 (n_136, n_110, n_111);
  xor g378 (n_469, n_112, n_113);
  xor g379 (n_119, n_469, in_2[8]);
  nand g380 (n_470, n_112, n_113);
  nand g381 (n_471, in_2[8], n_113);
  nand g382 (n_472, n_112, in_2[8]);
  nand g383 (n_139, n_470, n_471, n_472);
  xor g384 (n_473, in_3[8], n_116);
  xor g385 (n_123, n_473, n_117);
  nand g386 (n_474, in_3[8], n_116);
  nand g387 (n_475, n_117, n_116);
  nand g388 (n_476, in_3[8], n_117);
  nand g389 (n_142, n_474, n_475, n_476);
  xor g390 (n_477, n_118, n_119);
  xor g391 (n_126, n_477, n_120);
  nand g392 (n_478, n_118, n_119);
  nand g393 (n_479, n_120, n_119);
  nand g394 (n_480, n_118, n_120);
  nand g395 (n_145, n_478, n_479, n_480);
  xor g396 (n_481, n_121, n_122);
  xor g397 (n_129, n_481, n_123);
  nand g398 (n_482, n_121, n_122);
  nand g399 (n_483, n_123, n_122);
  nand g400 (n_484, n_121, n_123);
  nand g401 (n_148, n_482, n_483, n_484);
  xor g402 (n_485, n_124, n_125);
  xor g403 (n_131, n_485, n_126);
  nand g404 (n_486, n_124, n_125);
  nand g405 (n_487, n_126, n_125);
  nand g406 (n_488, n_124, n_126);
  nand g407 (n_152, n_486, n_487, n_488);
  xor g408 (n_489, n_127, n_128);
  xor g409 (n_132, n_489, n_129);
  nand g410 (n_490, n_127, n_128);
  nand g411 (n_491, n_129, n_128);
  nand g412 (n_492, n_127, n_129);
  nand g413 (n_154, n_490, n_491, n_492);
  xor g414 (n_493, n_130, n_131);
  xor g415 (out_1[8], n_493, n_132);
  nand g416 (n_494, n_130, n_131);
  nand g417 (n_495, n_132, n_131);
  nand g418 (n_496, n_130, n_132);
  nand g419 (out_0[9], n_494, n_495, n_496);
  xor g420 (n_497, n_133, in_2[9]);
  xor g421 (n_140, n_497, n_135);
  nand g422 (n_498, n_133, in_2[9]);
  nand g423 (n_499, n_135, in_2[9]);
  nand g424 (n_500, n_133, n_135);
  nand g425 (n_161, n_498, n_499, n_500);
  xor g426 (n_501, n_136, in_3[9]);
  xor g427 (n_144, n_501, n_138);
  nand g428 (n_502, n_136, in_3[9]);
  nand g429 (n_503, n_138, in_3[9]);
  nand g430 (n_504, n_136, n_138);
  nand g431 (n_164, n_502, n_503, n_504);
  xor g432 (n_505, n_139, n_140);
  xor g433 (n_146, n_505, n_141);
  nand g434 (n_506, n_139, n_140);
  nand g435 (n_507, n_141, n_140);
  nand g436 (n_508, n_139, n_141);
  nand g437 (n_166, n_506, n_507, n_508);
  xor g438 (n_509, n_142, n_143);
  xor g439 (n_151, n_509, n_144);
  nand g440 (n_510, n_142, n_143);
  nand g441 (n_511, n_144, n_143);
  nand g442 (n_512, n_142, n_144);
  nand g443 (n_169, n_510, n_511, n_512);
  xor g444 (n_513, n_145, n_146);
  xor g445 (n_153, n_513, n_147);
  nand g446 (n_514, n_145, n_146);
  nand g447 (n_515, n_147, n_146);
  nand g448 (n_516, n_145, n_147);
  nand g449 (n_174, n_514, n_515, n_516);
  xor g450 (n_517, n_148, n_149);
  xor g451 (n_155, n_517, n_150);
  nand g452 (n_518, n_148, n_149);
  nand g453 (n_519, n_150, n_149);
  nand g454 (n_520, n_148, n_150);
  nand g455 (n_177, n_518, n_519, n_520);
  xor g456 (n_521, n_151, n_152);
  xor g457 (n_156, n_521, n_153);
  nand g458 (n_522, n_151, n_152);
  nand g459 (n_523, n_153, n_152);
  nand g460 (n_524, n_151, n_153);
  nand g461 (n_178, n_522, n_523, n_524);
  xor g462 (n_525, n_154, n_155);
  xor g463 (out_1[9], n_525, n_156);
  nand g464 (n_526, n_154, n_155);
  nand g465 (n_527, n_156, n_155);
  nand g466 (n_528, n_154, n_156);
  nand g467 (out_0[10], n_526, n_527, n_528);
  xor g468 (n_529, n_157, in_2[10]);
  xor g469 (n_162, n_529, in_3[10]);
  nand g470 (n_530, n_157, in_2[10]);
  nand g471 (n_531, in_3[10], in_2[10]);
  nand g472 (n_532, n_157, in_3[10]);
  nand g473 (n_185, n_530, n_531, n_532);
  xor g474 (n_533, n_160, n_161);
  xor g475 (n_168, n_533, n_162);
  nand g476 (n_534, n_160, n_161);
  nand g477 (n_535, n_162, n_161);
  nand g478 (n_536, n_160, n_162);
  nand g479 (n_188, n_534, n_535, n_536);
  xor g480 (n_537, n_163, n_164);
  xor g481 (n_171, n_537, n_165);
  nand g482 (n_538, n_163, n_164);
  nand g483 (n_539, n_165, n_164);
  nand g484 (n_540, n_163, n_165);
  nand g485 (n_190, n_538, n_539, n_540);
  xor g486 (n_541, n_166, n_167);
  xor g487 (n_175, n_541, n_168);
  nand g488 (n_542, n_166, n_167);
  nand g489 (n_543, n_168, n_167);
  nand g490 (n_544, n_166, n_168);
  nand g491 (n_195, n_542, n_543, n_544);
  xor g492 (n_545, n_169, n_170);
  xor g493 (n_176, n_545, n_171);
  nand g494 (n_546, n_169, n_170);
  nand g495 (n_547, n_171, n_170);
  nand g496 (n_548, n_169, n_171);
  nand g497 (n_198, n_546, n_547, n_548);
  xor g498 (n_549, n_172, n_173);
  xor g499 (n_179, n_549, n_174);
  nand g500 (n_550, n_172, n_173);
  nand g501 (n_551, n_174, n_173);
  nand g502 (n_552, n_172, n_174);
  nand g503 (n_200, n_550, n_551, n_552);
  xor g504 (n_553, n_175, n_176);
  xor g505 (n_180, n_553, n_177);
  nand g506 (n_554, n_175, n_176);
  nand g507 (n_555, n_177, n_176);
  nand g508 (n_556, n_175, n_177);
  nand g509 (n_203, n_554, n_555, n_556);
  xor g510 (n_557, n_178, n_179);
  xor g511 (out_1[10], n_557, n_180);
  nand g512 (n_558, n_178, n_179);
  nand g513 (n_559, n_180, n_179);
  nand g514 (n_560, n_178, n_180);
  nand g515 (out_0[11], n_558, n_559, n_560);
  xor g516 (n_561, in_2[11], in_3[11]);
  xor g517 (n_186, n_561, n_183);
  nand g518 (n_562, in_2[11], in_3[11]);
  nand g519 (n_563, n_183, in_3[11]);
  nand g520 (n_564, in_2[11], n_183);
  nand g521 (n_209, n_562, n_563, n_564);
  xor g522 (n_565, n_184, n_185);
  xor g523 (n_192, n_565, n_186);
  nand g524 (n_566, n_184, n_185);
  nand g525 (n_567, n_186, n_185);
  nand g526 (n_568, n_184, n_186);
  nand g527 (n_212, n_566, n_567, n_568);
  xor g528 (n_569, n_187, n_188);
  xor g529 (n_197, n_569, n_189);
  nand g530 (n_570, n_187, n_188);
  nand g531 (n_571, n_189, n_188);
  nand g532 (n_572, n_187, n_189);
  nand g533 (n_216, n_570, n_571, n_572);
  xor g534 (n_573, n_190, n_191);
  xor g535 (n_199, n_573, n_192);
  nand g536 (n_574, n_190, n_191);
  nand g537 (n_575, n_192, n_191);
  nand g538 (n_576, n_190, n_192);
  nand g539 (n_218, n_574, n_575, n_576);
  xor g540 (n_577, n_193, n_194);
  xor g541 (n_201, n_577, n_195);
  nand g542 (n_578, n_193, n_194);
  nand g543 (n_579, n_195, n_194);
  nand g544 (n_580, n_193, n_195);
  nand g545 (n_222, n_578, n_579, n_580);
  xor g546 (n_581, n_196, n_197);
  xor g547 (n_202, n_581, n_198);
  nand g548 (n_582, n_196, n_197);
  nand g549 (n_583, n_198, n_197);
  nand g550 (n_584, n_196, n_198);
  nand g551 (n_225, n_582, n_583, n_584);
  xor g552 (n_585, n_199, n_200);
  xor g553 (n_204, n_585, n_201);
  nand g554 (n_586, n_199, n_200);
  nand g555 (n_587, n_201, n_200);
  nand g556 (n_588, n_199, n_201);
  nand g557 (n_227, n_586, n_587, n_588);
  xor g558 (n_589, n_202, n_203);
  xor g559 (out_1[11], n_589, n_204);
  nand g560 (n_590, n_202, n_203);
  nand g561 (n_591, n_204, n_203);
  nand g562 (n_592, n_202, n_204);
  nand g563 (out_0[12], n_590, n_591, n_592);
  xor g564 (n_593, in_2[12], in_3[12]);
  xor g565 (n_210, n_593, n_207);
  nand g566 (n_594, in_2[12], in_3[12]);
  nand g567 (n_595, n_207, in_3[12]);
  nand g568 (n_596, in_2[12], n_207);
  nand g569 (n_233, n_594, n_595, n_596);
  xor g570 (n_597, n_208, n_209);
  xor g571 (n_217, n_597, n_210);
  nand g572 (n_598, n_208, n_209);
  nand g573 (n_599, n_210, n_209);
  nand g574 (n_600, n_208, n_210);
  nand g575 (n_237, n_598, n_599, n_600);
  xor g576 (n_601, n_211, n_212);
  xor g577 (n_221, n_601, n_213);
  nand g578 (n_602, n_211, n_212);
  nand g579 (n_603, n_213, n_212);
  nand g580 (n_604, n_211, n_213);
  nand g581 (n_240, n_602, n_603, n_604);
  xor g582 (n_605, n_214, n_215);
  xor g583 (n_223, n_605, n_216);
  nand g584 (n_606, n_214, n_215);
  nand g585 (n_607, n_216, n_215);
  nand g586 (n_608, n_214, n_216);
  nand g587 (n_243, n_606, n_607, n_608);
  xor g588 (n_609, n_217, n_218);
  xor g589 (n_224, n_609, n_219);
  nand g590 (n_610, n_217, n_218);
  nand g591 (n_611, n_219, n_218);
  nand g592 (n_612, n_217, n_219);
  nand g593 (n_246, n_610, n_611, n_612);
  xor g594 (n_613, n_220, n_221);
  xor g595 (n_226, n_613, n_222);
  nand g596 (n_614, n_220, n_221);
  nand g597 (n_615, n_222, n_221);
  nand g598 (n_616, n_220, n_222);
  nand g599 (n_249, n_614, n_615, n_616);
  xor g600 (n_617, n_223, n_224);
  xor g601 (n_228, n_617, n_225);
  nand g602 (n_618, n_223, n_224);
  nand g603 (n_619, n_225, n_224);
  nand g604 (n_620, n_223, n_225);
  nand g605 (n_251, n_618, n_619, n_620);
  xor g606 (n_621, n_226, n_227);
  xor g607 (out_1[12], n_621, n_228);
  nand g608 (n_622, n_226, n_227);
  nand g609 (n_623, n_228, n_227);
  nand g610 (n_624, n_226, n_228);
  nand g611 (out_0[13], n_622, n_623, n_624);
  xor g612 (n_625, in_2[13], in_3[13]);
  xor g613 (n_234, n_625, n_231);
  nand g614 (n_626, in_2[13], in_3[13]);
  nand g615 (n_627, n_231, in_3[13]);
  nand g616 (n_628, in_2[13], n_231);
  nand g617 (n_257, n_626, n_627, n_628);
  xor g618 (n_629, n_232, n_233);
  xor g619 (n_241, n_629, n_234);
  nand g620 (n_630, n_232, n_233);
  nand g621 (n_631, n_234, n_233);
  nand g622 (n_632, n_232, n_234);
  nand g623 (n_261, n_630, n_631, n_632);
  xor g624 (n_633, n_235, n_236);
  xor g625 (n_244, n_633, n_237);
  nand g626 (n_634, n_235, n_236);
  nand g627 (n_635, n_237, n_236);
  nand g628 (n_636, n_235, n_237);
  nand g629 (n_265, n_634, n_635, n_636);
  xor g630 (n_637, n_238, n_239);
  xor g631 (n_247, n_637, n_240);
  nand g632 (n_638, n_238, n_239);
  nand g633 (n_639, n_240, n_239);
  nand g634 (n_640, n_238, n_240);
  nand g635 (n_269, n_638, n_639, n_640);
  xor g636 (n_641, n_241, n_242);
  xor g637 (n_248, n_641, n_243);
  nand g638 (n_642, n_241, n_242);
  nand g639 (n_643, n_243, n_242);
  nand g640 (n_644, n_241, n_243);
  nand g641 (n_270, n_642, n_643, n_644);
  xor g642 (n_645, n_244, n_245);
  xor g643 (n_250, n_645, n_246);
  nand g644 (n_646, n_244, n_245);
  nand g645 (n_647, n_246, n_245);
  nand g646 (n_648, n_244, n_246);
  nand g647 (n_272, n_646, n_647, n_648);
  xor g648 (n_649, n_247, n_248);
  xor g649 (n_252, n_649, n_249);
  nand g650 (n_650, n_247, n_248);
  nand g651 (n_651, n_249, n_248);
  nand g652 (n_652, n_247, n_249);
  nand g653 (n_274, n_650, n_651, n_652);
  xor g654 (n_653, n_250, n_251);
  xor g655 (out_1[13], n_653, n_252);
  nand g656 (n_654, n_250, n_251);
  nand g657 (n_655, n_252, n_251);
  nand g658 (n_656, n_250, n_252);
  nand g659 (out_0[14], n_654, n_655, n_656);
  xor g660 (n_657, in_2[14], in_3[14]);
  xor g661 (n_259, n_657, n_255);
  nand g662 (n_658, in_2[14], in_3[14]);
  nand g663 (n_659, n_255, in_3[14]);
  nand g664 (n_660, in_2[14], n_255);
  nand g665 (n_282, n_658, n_659, n_660);
  xor g666 (n_661, n_256, n_257);
  xor g667 (n_264, n_661, n_258);
  nand g668 (n_662, n_256, n_257);
  nand g669 (n_663, n_258, n_257);
  nand g670 (n_664, n_256, n_258);
  nand g671 (n_285, n_662, n_663, n_664);
  xor g672 (n_665, n_259, n_260);
  xor g673 (n_268, n_665, n_261);
  nand g674 (n_666, n_259, n_260);
  nand g675 (n_667, n_261, n_260);
  nand g676 (n_668, n_259, n_261);
  nand g677 (n_290, n_666, n_667, n_668);
  xor g678 (n_669, n_262, n_263);
  xor g679 (n_271, n_669, n_264);
  nand g680 (n_670, n_262, n_263);
  nand g681 (n_671, n_264, n_263);
  nand g682 (n_672, n_262, n_264);
  nand g683 (n_292, n_670, n_671, n_672);
  xor g684 (n_673, n_265, n_266);
  xor g685 (n_273, n_673, n_267);
  nand g686 (n_674, n_265, n_266);
  nand g687 (n_675, n_267, n_266);
  nand g688 (n_676, n_265, n_267);
  nand g689 (n_294, n_674, n_675, n_676);
  xor g690 (n_677, n_268, n_269);
  xor g691 (n_275, n_677, n_270);
  nand g692 (n_678, n_268, n_269);
  nand g693 (n_679, n_270, n_269);
  nand g694 (n_680, n_268, n_270);
  nand g695 (n_297, n_678, n_679, n_680);
  xor g696 (n_681, n_271, n_272);
  xor g697 (n_276, n_681, n_273);
  nand g698 (n_682, n_271, n_272);
  nand g699 (n_683, n_273, n_272);
  nand g700 (n_684, n_271, n_273);
  nand g701 (n_299, n_682, n_683, n_684);
  xor g702 (n_685, n_274, n_275);
  xor g703 (out_1[14], n_685, n_276);
  nand g704 (n_686, n_274, n_275);
  nand g705 (n_687, n_276, n_275);
  nand g706 (n_688, n_274, n_276);
  nand g707 (out_0[15], n_686, n_687, n_688);
  xor g708 (n_689, in_2[15], in_3[15]);
  xor g709 (n_283, n_689, n_279);
  nand g710 (n_690, in_2[15], in_3[15]);
  nand g711 (n_691, n_279, in_3[15]);
  nand g712 (n_692, in_2[15], n_279);
  nand g713 (n_303, n_690, n_691, n_692);
  xor g714 (n_693, n_280, n_281);
  xor g715 (n_291, n_693, n_282);
  nand g716 (n_694, n_280, n_281);
  nand g717 (n_695, n_282, n_281);
  nand g718 (n_696, n_280, n_282);
  nand g719 (n_308, n_694, n_695, n_696);
  xor g720 (n_697, n_283, n_284);
  xor g721 (n_293, n_697, n_285);
  nand g722 (n_698, n_283, n_284);
  nand g723 (n_699, n_285, n_284);
  nand g724 (n_700, n_283, n_285);
  nand g725 (n_311, n_698, n_699, n_700);
  xor g726 (n_701, n_286, n_287);
  xor g727 (n_295, n_701, n_288);
  nand g728 (n_702, n_286, n_287);
  nand g729 (n_703, n_288, n_287);
  nand g730 (n_704, n_286, n_288);
  nand g731 (n_312, n_702, n_703, n_704);
  xor g732 (n_705, n_289, n_290);
  xor g733 (n_296, n_705, n_291);
  nand g734 (n_706, n_289, n_290);
  nand g735 (n_707, n_291, n_290);
  nand g736 (n_708, n_289, n_291);
  nand g737 (n_315, n_706, n_707, n_708);
  xor g738 (n_709, n_292, n_293);
  xor g739 (n_298, n_709, n_294);
  nand g740 (n_710, n_292, n_293);
  nand g741 (n_711, n_294, n_293);
  nand g742 (n_712, n_292, n_294);
  nand g743 (n_318, n_710, n_711, n_712);
  xor g744 (n_713, n_295, n_296);
  xor g745 (n_300, n_713, n_297);
  nand g746 (n_714, n_295, n_296);
  nand g747 (n_715, n_297, n_296);
  nand g748 (n_716, n_295, n_297);
  nand g749 (n_320, n_714, n_715, n_716);
  xor g750 (n_717, n_298, n_299);
  xor g751 (out_1[15], n_717, n_300);
  nand g752 (n_718, n_298, n_299);
  nand g753 (n_719, n_300, n_299);
  nand g754 (n_720, n_298, n_300);
  nand g755 (out_0[16], n_718, n_719, n_720);
  xor g756 (n_721, n_301, n_302);
  xor g757 (n_309, n_721, n_303);
  xor g762 (n_725, n_304, n_305);
  xor g763 (n_313, n_725, n_306);
  xor g768 (n_729, n_307, n_308);
  xor g769 (n_316, n_729, n_309);
  xor g774 (n_733, n_310, n_311);
  xor g775 (n_317, n_733, n_312);
  xor g780 (n_737, n_313, n_314);
  xor g781 (n_319, n_737, n_315);
  xor g786 (n_741, n_316, n_317);
  xor g787 (n_321, n_741, n_318);
  xor g792 (n_745, n_319, n_320);
  xor g793 (out_1[16], n_745, n_321);
endmodule

module csa_tree_271_GENERIC(in_0, in_1, in_2, in_3, out_0, out_1,
     out_2);
  input [16:0] in_0, in_2, in_3;
  input [7:0] in_1;
  output [16:0] out_0, out_1;
  output out_2;
  wire [16:0] in_0, in_2, in_3;
  wire [7:0] in_1;
  wire [16:0] out_0, out_1;
  wire out_2;
  csa_tree_271_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .in_3 (in_3), .out_0 (out_0), .out_1 (out_1), .out_2
       (out_2));
endmodule

module csa_tree_mul_25_40_group_52_GENERIC_REAL(in_0, in_1, out_0);
// synthesis_equation "assign out_0 = ( in_0 * in_1 )  ;"
  input [15:0] in_0;
  input [7:0] in_1;
  output [16:0] out_0;
  wire [15:0] in_0;
  wire [7:0] in_1;
  wire [16:0] out_0;
  wire n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
  wire n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187;
  wire n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195;
  wire n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203;
  wire n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211;
  wire n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219;
  wire n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227;
  wire n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251;
  wire n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259;
  wire n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267;
  wire n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275;
  wire n_276, n_277, n_278, n_279, n_280, n_281, n_282, n_283;
  wire n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291;
  wire n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299;
  wire n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307;
  wire n_308, n_309, n_310, n_311, n_312, n_313, n_314, n_315;
  wire n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323;
  wire n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339;
  wire n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347;
  wire n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
  wire n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459;
  wire n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475;
  wire n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483;
  wire n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491;
  wire n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499;
  wire n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515;
  wire n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523;
  wire n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_550;
  wire n_554, n_558, n_562, n_569, n_572, n_574, n_577, n_579;
  wire n_580, n_582, n_584, n_585, n_587, n_589, n_590, n_592;
  wire n_594, n_595, n_597, n_599, n_600, n_602, n_604, n_605;
  wire n_607, n_609, n_610, n_612, n_614, n_615, n_617, n_619;
  wire n_620, n_622, n_624, n_625, n_627, n_629, n_630, n_632;
  wire n_634, n_635, n_637, n_639, n_640, n_642, n_644, n_645;
  wire n_647, n_668, n_670, n_671, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  and g1 (out_0[0], in_0[0], in_1[0]);
  and g2 (n_57, in_0[1], in_1[0]);
  and g3 (n_77, in_0[2], in_1[0]);
  and g4 (n_79, in_0[3], in_1[0]);
  and g5 (n_84, in_0[4], in_1[0]);
  and g6 (n_92, in_0[5], in_1[0]);
  and g7 (n_103, in_0[6], in_1[0]);
  and g8 (n_117, in_0[7], in_1[0]);
  and g9 (n_133, in_0[8], in_1[0]);
  and g10 (n_151, in_0[9], in_1[0]);
  and g11 (n_169, in_0[10], in_1[0]);
  and g12 (n_187, in_0[11], in_1[0]);
  and g13 (n_205, in_0[12], in_1[0]);
  and g14 (n_223, in_0[13], in_1[0]);
  and g15 (n_241, in_0[14], in_1[0]);
  and g16 (n_259, in_0[15], in_1[0]);
  and g17 (n_74, in_0[0], in_1[1]);
  and g18 (n_56, in_0[1], in_1[1]);
  and g19 (n_80, in_0[2], in_1[1]);
  and g20 (n_85, in_0[3], in_1[1]);
  and g21 (n_93, in_0[4], in_1[1]);
  and g22 (n_104, in_0[5], in_1[1]);
  and g23 (n_118, in_0[6], in_1[1]);
  and g24 (n_134, in_0[7], in_1[1]);
  and g25 (n_152, in_0[8], in_1[1]);
  and g26 (n_170, in_0[9], in_1[1]);
  and g27 (n_188, in_0[10], in_1[1]);
  and g28 (n_206, in_0[11], in_1[1]);
  and g29 (n_224, in_0[12], in_1[1]);
  and g30 (n_242, in_0[13], in_1[1]);
  and g31 (n_260, in_0[14], in_1[1]);
  and g32 (n_277, in_0[15], in_1[1]);
  and g33 (n_78, in_0[0], in_1[2]);
  and g34 (n_82, in_0[1], in_1[2]);
  and g35 (n_88, in_0[2], in_1[2]);
  and g36 (n_96, in_0[3], in_1[2]);
  and g37 (n_107, in_0[4], in_1[2]);
  and g38 (n_122, in_0[5], in_1[2]);
  and g39 (n_138, in_0[6], in_1[2]);
  and g40 (n_156, in_0[7], in_1[2]);
  and g41 (n_174, in_0[8], in_1[2]);
  and g42 (n_192, in_0[9], in_1[2]);
  and g43 (n_210, in_0[10], in_1[2]);
  and g44 (n_228, in_0[11], in_1[2]);
  and g45 (n_246, in_0[12], in_1[2]);
  and g46 (n_264, in_0[13], in_1[2]);
  and g47 (n_278, in_0[14], in_1[2]);
  and g48 (n_81, in_0[0], in_1[3]);
  and g49 (n_86, in_0[1], in_1[3]);
  and g50 (n_94, in_0[2], in_1[3]);
  and g51 (n_105, in_0[3], in_1[3]);
  and g52 (n_119, in_0[4], in_1[3]);
  and g53 (n_135, in_0[5], in_1[3]);
  and g54 (n_153, in_0[6], in_1[3]);
  and g55 (n_171, in_0[7], in_1[3]);
  and g56 (n_189, in_0[8], in_1[3]);
  and g57 (n_207, in_0[9], in_1[3]);
  and g58 (n_225, in_0[10], in_1[3]);
  and g59 (n_243, in_0[11], in_1[3]);
  and g60 (n_261, in_0[12], in_1[3]);
  and g61 (n_281, in_0[13], in_1[3]);
  and g62 (n_87, in_0[0], in_1[4]);
  and g63 (n_95, in_0[1], in_1[4]);
  and g64 (n_106, in_0[2], in_1[4]);
  and g65 (n_121, in_0[3], in_1[4]);
  and g66 (n_137, in_0[4], in_1[4]);
  and g67 (n_155, in_0[5], in_1[4]);
  and g68 (n_173, in_0[6], in_1[4]);
  and g69 (n_191, in_0[7], in_1[4]);
  and g70 (n_209, in_0[8], in_1[4]);
  and g71 (n_227, in_0[9], in_1[4]);
  and g72 (n_245, in_0[10], in_1[4]);
  and g73 (n_263, in_0[11], in_1[4]);
  and g74 (n_279, in_0[12], in_1[4]);
  and g75 (n_97, in_0[0], in_1[5]);
  and g76 (n_108, in_0[1], in_1[5]);
  and g77 (n_123, in_0[2], in_1[5]);
  and g78 (n_139, in_0[3], in_1[5]);
  and g79 (n_157, in_0[4], in_1[5]);
  and g80 (n_175, in_0[5], in_1[5]);
  and g81 (n_193, in_0[6], in_1[5]);
  and g82 (n_211, in_0[7], in_1[5]);
  and g83 (n_229, in_0[8], in_1[5]);
  and g84 (n_247, in_0[9], in_1[5]);
  and g85 (n_265, in_0[10], in_1[5]);
  and g86 (n_280, in_0[11], in_1[5]);
  and g87 (n_109, in_0[0], in_1[6]);
  and g88 (n_124, in_0[1], in_1[6]);
  and g89 (n_140, in_0[2], in_1[6]);
  and g90 (n_158, in_0[3], in_1[6]);
  and g91 (n_176, in_0[4], in_1[6]);
  and g92 (n_194, in_0[5], in_1[6]);
  and g93 (n_212, in_0[6], in_1[6]);
  and g94 (n_230, in_0[7], in_1[6]);
  and g95 (n_248, in_0[8], in_1[6]);
  and g96 (n_266, in_0[9], in_1[6]);
  and g97 (n_282, in_0[10], in_1[6]);
  and g98 (n_120, in_0[0], in_1[7]);
  and g99 (n_136, in_0[1], in_1[7]);
  and g100 (n_154, in_0[2], in_1[7]);
  and g101 (n_172, in_0[3], in_1[7]);
  and g102 (n_190, in_0[4], in_1[7]);
  and g103 (n_208, in_0[5], in_1[7]);
  and g104 (n_226, in_0[6], in_1[7]);
  and g105 (n_244, in_0[7], in_1[7]);
  and g106 (n_262, in_0[8], in_1[7]);
  and g107 (n_283, in_0[9], in_1[7]);
  xor g183 (n_73, n_77, n_78);
  and g184 (n_55, n_77, n_78);
  xor g185 (n_83, n_79, n_80);
  and g186 (n_90, n_79, n_80);
  xor g187 (n_294, n_81, n_82);
  xor g188 (n_72, n_294, n_83);
  nand g189 (n_295, n_81, n_82);
  nand g190 (n_296, n_83, n_82);
  nand g191 (n_297, n_81, n_83);
  nand g192 (n_54, n_295, n_296, n_297);
  xor g193 (n_89, n_84, n_85);
  and g194 (n_99, n_84, n_85);
  xor g195 (n_298, n_86, n_87);
  xor g196 (n_91, n_298, n_88);
  nand g197 (n_299, n_86, n_87);
  nand g198 (n_300, n_88, n_87);
  nand g199 (n_301, n_86, n_88);
  nand g200 (n_100, n_299, n_300, n_301);
  xor g201 (n_302, n_89, n_90);
  xor g202 (n_71, n_302, n_91);
  nand g203 (n_303, n_89, n_90);
  nand g204 (n_304, n_91, n_90);
  nand g205 (n_305, n_89, n_91);
  nand g206 (n_53, n_303, n_304, n_305);
  xor g207 (n_98, n_92, n_93);
  and g208 (n_110, n_92, n_93);
  xor g209 (n_306, n_94, n_95);
  xor g210 (n_101, n_306, n_96);
  nand g211 (n_307, n_94, n_95);
  nand g212 (n_308, n_96, n_95);
  nand g213 (n_309, n_94, n_96);
  nand g214 (n_112, n_307, n_308, n_309);
  xor g215 (n_310, n_97, n_98);
  xor g216 (n_102, n_310, n_99);
  nand g217 (n_311, n_97, n_98);
  nand g218 (n_312, n_99, n_98);
  nand g219 (n_313, n_97, n_99);
  nand g220 (n_114, n_311, n_312, n_313);
  xor g221 (n_314, n_100, n_101);
  xor g222 (n_70, n_314, n_102);
  nand g223 (n_315, n_100, n_101);
  nand g224 (n_316, n_102, n_101);
  nand g225 (n_317, n_100, n_102);
  nand g226 (n_52, n_315, n_316, n_317);
  xor g227 (n_111, n_103, n_104);
  and g228 (n_125, n_103, n_104);
  xor g229 (n_318, n_105, n_106);
  xor g230 (n_113, n_318, n_107);
  nand g231 (n_319, n_105, n_106);
  nand g232 (n_320, n_107, n_106);
  nand g233 (n_321, n_105, n_107);
  nand g234 (n_75, n_319, n_320, n_321);
  xor g235 (n_322, n_108, n_109);
  xor g236 (n_115, n_322, n_110);
  nand g237 (n_323, n_108, n_109);
  nand g238 (n_324, n_110, n_109);
  nand g239 (n_325, n_108, n_110);
  nand g240 (n_129, n_323, n_324, n_325);
  xor g241 (n_326, n_111, n_112);
  xor g242 (n_116, n_326, n_113);
  nand g243 (n_327, n_111, n_112);
  nand g244 (n_328, n_113, n_112);
  nand g245 (n_329, n_111, n_113);
  nand g246 (n_131, n_327, n_328, n_329);
  xor g247 (n_330, n_114, n_115);
  xor g248 (n_69, n_330, n_116);
  nand g249 (n_331, n_114, n_115);
  nand g250 (n_332, n_116, n_115);
  nand g251 (n_333, n_114, n_116);
  nand g252 (n_51, n_331, n_332, n_333);
  xor g253 (n_126, n_117, n_118);
  and g254 (n_141, n_117, n_118);
  xor g255 (n_334, n_119, n_120);
  xor g256 (n_128, n_334, n_121);
  nand g257 (n_335, n_119, n_120);
  nand g258 (n_336, n_121, n_120);
  nand g259 (n_337, n_119, n_121);
  nand g260 (n_142, n_335, n_336, n_337);
  xor g261 (n_338, n_122, n_123);
  xor g262 (n_127, n_338, n_124);
  nand g263 (n_339, n_122, n_123);
  nand g264 (n_340, n_124, n_123);
  nand g265 (n_341, n_122, n_124);
  nand g266 (n_143, n_339, n_340, n_341);
  xor g267 (n_342, n_125, n_126);
  xor g268 (n_130, n_342, n_75);
  nand g269 (n_343, n_125, n_126);
  nand g270 (n_344, n_75, n_126);
  nand g271 (n_345, n_125, n_75);
  nand g272 (n_147, n_343, n_344, n_345);
  xor g273 (n_346, n_127, n_128);
  xor g274 (n_132, n_346, n_129);
  nand g275 (n_347, n_127, n_128);
  nand g276 (n_348, n_129, n_128);
  nand g277 (n_349, n_127, n_129);
  nand g278 (n_149, n_347, n_348, n_349);
  xor g279 (n_350, n_130, n_131);
  xor g280 (n_68, n_350, n_132);
  nand g281 (n_351, n_130, n_131);
  nand g282 (n_352, n_132, n_131);
  nand g283 (n_353, n_130, n_132);
  nand g284 (n_50, n_351, n_352, n_353);
  xor g285 (n_354, n_133, n_134);
  xor g286 (n_144, n_354, n_135);
  nand g287 (n_355, n_133, n_134);
  nand g288 (n_356, n_135, n_134);
  nand g289 (n_357, n_133, n_135);
  nand g290 (n_159, n_355, n_356, n_357);
  xor g291 (n_358, n_136, n_137);
  xor g292 (n_145, n_358, n_138);
  nand g293 (n_359, n_136, n_137);
  nand g294 (n_360, n_138, n_137);
  nand g295 (n_361, n_136, n_138);
  nand g296 (n_160, n_359, n_360, n_361);
  xor g297 (n_362, n_139, n_140);
  xor g298 (n_146, n_362, n_141);
  nand g299 (n_363, n_139, n_140);
  nand g300 (n_364, n_141, n_140);
  nand g301 (n_365, n_139, n_141);
  nand g302 (n_163, n_363, n_364, n_365);
  xor g303 (n_366, n_142, n_143);
  xor g304 (n_148, n_366, n_144);
  nand g305 (n_367, n_142, n_143);
  nand g306 (n_368, n_144, n_143);
  nand g307 (n_369, n_142, n_144);
  nand g308 (n_165, n_367, n_368, n_369);
  xor g309 (n_370, n_145, n_146);
  xor g310 (n_150, n_370, n_147);
  nand g311 (n_371, n_145, n_146);
  nand g312 (n_372, n_147, n_146);
  nand g313 (n_373, n_145, n_147);
  nand g314 (n_167, n_371, n_372, n_373);
  xor g315 (n_374, n_148, n_149);
  xor g316 (n_67, n_374, n_150);
  nand g317 (n_375, n_148, n_149);
  nand g318 (n_376, n_150, n_149);
  nand g319 (n_377, n_148, n_150);
  nand g320 (n_49, n_375, n_376, n_377);
  xor g321 (n_378, n_151, n_152);
  xor g322 (n_161, n_378, n_153);
  nand g323 (n_379, n_151, n_152);
  nand g324 (n_380, n_153, n_152);
  nand g325 (n_381, n_151, n_153);
  nand g326 (n_177, n_379, n_380, n_381);
  xor g327 (n_382, n_154, n_155);
  xor g328 (n_162, n_382, n_156);
  nand g329 (n_383, n_154, n_155);
  nand g330 (n_384, n_156, n_155);
  nand g331 (n_385, n_154, n_156);
  nand g332 (n_178, n_383, n_384, n_385);
  xor g333 (n_386, n_157, n_158);
  xor g334 (n_164, n_386, n_159);
  nand g335 (n_387, n_157, n_158);
  nand g336 (n_388, n_159, n_158);
  nand g337 (n_389, n_157, n_159);
  nand g338 (n_182, n_387, n_388, n_389);
  xor g339 (n_390, n_160, n_161);
  xor g340 (n_166, n_390, n_162);
  nand g341 (n_391, n_160, n_161);
  nand g342 (n_392, n_162, n_161);
  nand g343 (n_393, n_160, n_162);
  nand g344 (n_183, n_391, n_392, n_393);
  xor g345 (n_394, n_163, n_164);
  xor g346 (n_168, n_394, n_165);
  nand g347 (n_395, n_163, n_164);
  nand g348 (n_396, n_165, n_164);
  nand g349 (n_397, n_163, n_165);
  nand g350 (n_186, n_395, n_396, n_397);
  xor g351 (n_398, n_166, n_167);
  xor g352 (n_66, n_398, n_168);
  nand g353 (n_399, n_166, n_167);
  nand g354 (n_400, n_168, n_167);
  nand g355 (n_401, n_166, n_168);
  nand g356 (n_48, n_399, n_400, n_401);
  xor g357 (n_402, n_169, n_170);
  xor g358 (n_179, n_402, n_171);
  nand g359 (n_403, n_169, n_170);
  nand g360 (n_404, n_171, n_170);
  nand g361 (n_405, n_169, n_171);
  nand g362 (n_195, n_403, n_404, n_405);
  xor g363 (n_406, n_172, n_173);
  xor g364 (n_180, n_406, n_174);
  nand g365 (n_407, n_172, n_173);
  nand g366 (n_408, n_174, n_173);
  nand g367 (n_409, n_172, n_174);
  nand g368 (n_196, n_407, n_408, n_409);
  xor g369 (n_410, n_175, n_176);
  xor g370 (n_181, n_410, n_177);
  nand g371 (n_411, n_175, n_176);
  nand g372 (n_412, n_177, n_176);
  nand g373 (n_413, n_175, n_177);
  nand g374 (n_200, n_411, n_412, n_413);
  xor g375 (n_414, n_178, n_179);
  xor g376 (n_184, n_414, n_180);
  nand g377 (n_415, n_178, n_179);
  nand g378 (n_416, n_180, n_179);
  nand g379 (n_417, n_178, n_180);
  nand g380 (n_201, n_415, n_416, n_417);
  xor g381 (n_418, n_181, n_182);
  xor g382 (n_185, n_418, n_183);
  nand g383 (n_419, n_181, n_182);
  nand g384 (n_420, n_183, n_182);
  nand g385 (n_421, n_181, n_183);
  nand g386 (n_204, n_419, n_420, n_421);
  xor g387 (n_422, n_184, n_185);
  xor g388 (n_65, n_422, n_186);
  nand g389 (n_423, n_184, n_185);
  nand g390 (n_424, n_186, n_185);
  nand g391 (n_425, n_184, n_186);
  nand g392 (n_47, n_423, n_424, n_425);
  xor g393 (n_426, n_187, n_188);
  xor g394 (n_197, n_426, n_189);
  nand g395 (n_427, n_187, n_188);
  nand g396 (n_428, n_189, n_188);
  nand g397 (n_429, n_187, n_189);
  nand g398 (n_213, n_427, n_428, n_429);
  xor g399 (n_430, n_190, n_191);
  xor g400 (n_198, n_430, n_192);
  nand g401 (n_431, n_190, n_191);
  nand g402 (n_432, n_192, n_191);
  nand g403 (n_433, n_190, n_192);
  nand g404 (n_214, n_431, n_432, n_433);
  xor g405 (n_434, n_193, n_194);
  xor g406 (n_199, n_434, n_195);
  nand g407 (n_435, n_193, n_194);
  nand g408 (n_436, n_195, n_194);
  nand g409 (n_437, n_193, n_195);
  nand g410 (n_218, n_435, n_436, n_437);
  xor g411 (n_438, n_196, n_197);
  xor g412 (n_202, n_438, n_198);
  nand g413 (n_439, n_196, n_197);
  nand g414 (n_440, n_198, n_197);
  nand g415 (n_441, n_196, n_198);
  nand g416 (n_219, n_439, n_440, n_441);
  xor g417 (n_442, n_199, n_200);
  xor g418 (n_203, n_442, n_201);
  nand g419 (n_443, n_199, n_200);
  nand g420 (n_444, n_201, n_200);
  nand g421 (n_445, n_199, n_201);
  nand g422 (n_222, n_443, n_444, n_445);
  xor g423 (n_446, n_202, n_203);
  xor g424 (n_64, n_446, n_204);
  nand g425 (n_447, n_202, n_203);
  nand g426 (n_448, n_204, n_203);
  nand g427 (n_449, n_202, n_204);
  nand g428 (n_46, n_447, n_448, n_449);
  xor g429 (n_450, n_205, n_206);
  xor g430 (n_215, n_450, n_207);
  nand g431 (n_451, n_205, n_206);
  nand g432 (n_452, n_207, n_206);
  nand g433 (n_453, n_205, n_207);
  nand g434 (n_231, n_451, n_452, n_453);
  xor g435 (n_454, n_208, n_209);
  xor g436 (n_216, n_454, n_210);
  nand g437 (n_455, n_208, n_209);
  nand g438 (n_456, n_210, n_209);
  nand g439 (n_457, n_208, n_210);
  nand g440 (n_232, n_455, n_456, n_457);
  xor g441 (n_458, n_211, n_212);
  xor g442 (n_217, n_458, n_213);
  nand g443 (n_459, n_211, n_212);
  nand g444 (n_460, n_213, n_212);
  nand g445 (n_461, n_211, n_213);
  nand g446 (n_236, n_459, n_460, n_461);
  xor g447 (n_462, n_214, n_215);
  xor g448 (n_220, n_462, n_216);
  nand g449 (n_463, n_214, n_215);
  nand g450 (n_464, n_216, n_215);
  nand g451 (n_465, n_214, n_216);
  nand g452 (n_237, n_463, n_464, n_465);
  xor g453 (n_466, n_217, n_218);
  xor g454 (n_221, n_466, n_219);
  nand g455 (n_467, n_217, n_218);
  nand g456 (n_468, n_219, n_218);
  nand g457 (n_469, n_217, n_219);
  nand g458 (n_240, n_467, n_468, n_469);
  xor g459 (n_470, n_220, n_221);
  xor g460 (n_63, n_470, n_222);
  nand g461 (n_471, n_220, n_221);
  nand g462 (n_472, n_222, n_221);
  nand g463 (n_473, n_220, n_222);
  nand g464 (n_45, n_471, n_472, n_473);
  xor g465 (n_474, n_223, n_224);
  xor g466 (n_233, n_474, n_225);
  nand g467 (n_475, n_223, n_224);
  nand g468 (n_476, n_225, n_224);
  nand g469 (n_477, n_223, n_225);
  nand g470 (n_249, n_475, n_476, n_477);
  xor g471 (n_478, n_226, n_227);
  xor g472 (n_234, n_478, n_228);
  nand g473 (n_479, n_226, n_227);
  nand g474 (n_480, n_228, n_227);
  nand g475 (n_481, n_226, n_228);
  nand g476 (n_250, n_479, n_480, n_481);
  xor g477 (n_482, n_229, n_230);
  xor g478 (n_235, n_482, n_231);
  nand g479 (n_483, n_229, n_230);
  nand g480 (n_484, n_231, n_230);
  nand g481 (n_485, n_229, n_231);
  nand g482 (n_254, n_483, n_484, n_485);
  xor g483 (n_486, n_232, n_233);
  xor g484 (n_238, n_486, n_234);
  nand g485 (n_487, n_232, n_233);
  nand g486 (n_488, n_234, n_233);
  nand g487 (n_489, n_232, n_234);
  nand g488 (n_255, n_487, n_488, n_489);
  xor g489 (n_490, n_235, n_236);
  xor g490 (n_239, n_490, n_237);
  nand g491 (n_491, n_235, n_236);
  nand g492 (n_492, n_237, n_236);
  nand g493 (n_493, n_235, n_237);
  nand g494 (n_258, n_491, n_492, n_493);
  xor g495 (n_494, n_238, n_239);
  xor g496 (n_62, n_494, n_240);
  nand g497 (n_495, n_238, n_239);
  nand g498 (n_496, n_240, n_239);
  nand g499 (n_497, n_238, n_240);
  nand g500 (n_44, n_495, n_496, n_497);
  xor g501 (n_498, n_241, n_242);
  xor g502 (n_251, n_498, n_243);
  nand g503 (n_499, n_241, n_242);
  nand g504 (n_500, n_243, n_242);
  nand g505 (n_501, n_241, n_243);
  nand g506 (n_267, n_499, n_500, n_501);
  xor g507 (n_502, n_244, n_245);
  xor g508 (n_252, n_502, n_246);
  nand g509 (n_503, n_244, n_245);
  nand g510 (n_504, n_246, n_245);
  nand g511 (n_505, n_244, n_246);
  nand g512 (n_268, n_503, n_504, n_505);
  xor g513 (n_506, n_247, n_248);
  xor g514 (n_253, n_506, n_249);
  nand g515 (n_507, n_247, n_248);
  nand g516 (n_508, n_249, n_248);
  nand g517 (n_509, n_247, n_249);
  nand g518 (n_272, n_507, n_508, n_509);
  xor g519 (n_510, n_250, n_251);
  xor g520 (n_256, n_510, n_252);
  nand g521 (n_511, n_250, n_251);
  nand g522 (n_512, n_252, n_251);
  nand g523 (n_513, n_250, n_252);
  nand g524 (n_273, n_511, n_512, n_513);
  xor g525 (n_514, n_253, n_254);
  xor g526 (n_257, n_514, n_255);
  nand g527 (n_515, n_253, n_254);
  nand g528 (n_516, n_255, n_254);
  nand g529 (n_517, n_253, n_255);
  nand g530 (n_276, n_515, n_516, n_517);
  xor g531 (n_518, n_256, n_257);
  xor g532 (n_61, n_518, n_258);
  nand g533 (n_519, n_256, n_257);
  nand g534 (n_520, n_258, n_257);
  nand g535 (n_521, n_256, n_258);
  nand g536 (n_43, n_519, n_520, n_521);
  xor g537 (n_522, n_259, n_260);
  xor g538 (n_269, n_522, n_261);
  nand g539 (n_523, n_259, n_260);
  nand g540 (n_524, n_261, n_260);
  nand g541 (n_525, n_259, n_261);
  nand g542 (n_286, n_523, n_524, n_525);
  xor g543 (n_526, n_262, n_263);
  xor g544 (n_270, n_526, n_264);
  nand g545 (n_527, n_262, n_263);
  nand g546 (n_528, n_264, n_263);
  nand g547 (n_529, n_262, n_264);
  nand g548 (n_285, n_527, n_528, n_529);
  xor g549 (n_530, n_265, n_266);
  xor g550 (n_271, n_530, n_267);
  nand g551 (n_531, n_265, n_266);
  nand g552 (n_532, n_267, n_266);
  nand g553 (n_533, n_265, n_267);
  nand g554 (n_289, n_531, n_532, n_533);
  xor g555 (n_534, n_268, n_269);
  xor g556 (n_274, n_534, n_270);
  nand g557 (n_535, n_268, n_269);
  nand g558 (n_536, n_270, n_269);
  nand g559 (n_537, n_268, n_270);
  nand g560 (n_290, n_535, n_536, n_537);
  xor g561 (n_538, n_271, n_272);
  xor g562 (n_275, n_538, n_273);
  nand g563 (n_539, n_271, n_272);
  nand g564 (n_540, n_273, n_272);
  nand g565 (n_541, n_271, n_273);
  nand g566 (n_293, n_539, n_540, n_541);
  xor g567 (n_542, n_274, n_275);
  xor g568 (n_60, n_542, n_276);
  nand g569 (n_543, n_274, n_275);
  nand g570 (n_544, n_276, n_275);
  nand g571 (n_545, n_274, n_276);
  nand g572 (n_42, n_543, n_544, n_545);
  xor g573 (n_284, n_277, n_278);
  xor g575 (n_546, n_279, n_280);
  xor g576 (n_287, n_546, n_281);
  xor g581 (n_550, n_282, n_283);
  xor g582 (n_288, n_550, n_284);
  xor g587 (n_554, n_285, n_286);
  xor g588 (n_291, n_554, n_287);
  xor g593 (n_558, n_288, n_289);
  xor g594 (n_292, n_558, n_290);
  xor g599 (n_562, n_291, n_292);
  xor g600 (n_59, n_562, n_293);
  nor g610 (n_569, n_57, n_74);
  nand g611 (n_572, n_57, n_74);
  nor g612 (n_574, n_56, n_73);
  nand g613 (n_577, n_56, n_73);
  nor g614 (n_579, n_55, n_72);
  nand g615 (n_582, n_55, n_72);
  nor g616 (n_584, n_54, n_71);
  nand g617 (n_587, n_54, n_71);
  nor g618 (n_589, n_53, n_70);
  nand g619 (n_592, n_53, n_70);
  nor g620 (n_594, n_52, n_69);
  nand g621 (n_597, n_52, n_69);
  nor g622 (n_599, n_51, n_68);
  nand g623 (n_602, n_51, n_68);
  nor g624 (n_604, n_50, n_67);
  nand g625 (n_607, n_50, n_67);
  nor g626 (n_609, n_49, n_66);
  nand g627 (n_612, n_49, n_66);
  nor g628 (n_614, n_48, n_65);
  nand g629 (n_617, n_48, n_65);
  nor g630 (n_619, n_47, n_64);
  nand g631 (n_622, n_47, n_64);
  nor g632 (n_624, n_46, n_63);
  nand g633 (n_627, n_46, n_63);
  nor g634 (n_629, n_45, n_62);
  nand g635 (n_632, n_45, n_62);
  nor g636 (n_634, n_44, n_61);
  nand g637 (n_637, n_44, n_61);
  nor g638 (n_639, n_43, n_60);
  nand g639 (n_642, n_43, n_60);
  nor g640 (n_644, n_42, n_59);
  nand g641 (n_647, n_42, n_59);
  nand g647 (n_580, n_577, n_671);
  nand g650 (n_585, n_582, n_675);
  nand g653 (n_590, n_587, n_678);
  nand g656 (n_595, n_592, n_681);
  nand g659 (n_600, n_597, n_690);
  nand g662 (n_605, n_602, n_691);
  nand g665 (n_610, n_607, n_692);
  nand g668 (n_615, n_612, n_693);
  nand g671 (n_620, n_617, n_694);
  nand g674 (n_625, n_622, n_695);
  nand g677 (n_630, n_627, n_696);
  nand g680 (n_635, n_632, n_697);
  nand g683 (n_640, n_637, n_698);
  nand g686 (n_645, n_642, n_699);
  xnor g693 (out_0[3], n_580, n_673);
  xnor g695 (out_0[4], n_585, n_674);
  xnor g697 (out_0[5], n_590, n_676);
  xnor g699 (out_0[6], n_595, n_677);
  xnor g701 (out_0[7], n_600, n_679);
  xnor g703 (out_0[8], n_605, n_680);
  xnor g705 (out_0[9], n_610, n_682);
  xnor g707 (out_0[10], n_615, n_683);
  xnor g709 (out_0[11], n_620, n_684);
  xnor g109 (out_0[12], n_625, n_685);
  xnor g111 (out_0[13], n_630, n_686);
  xnor g113 (out_0[14], n_635, n_687);
  xnor g115 (out_0[15], n_640, n_688);
  xnor g117 (out_0[16], n_645, n_689);
  or g710 (n_668, wc, n_569);
  not gc (wc, n_572);
  not g712 (out_0[1], n_668);
  or g713 (n_670, wc0, n_574);
  not gc0 (wc0, n_577);
  or g714 (n_671, n_572, n_574);
  xor g715 (out_0[2], n_572, n_670);
  or g716 (n_673, wc1, n_579);
  not gc1 (wc1, n_582);
  or g717 (n_674, wc2, n_584);
  not gc2 (wc2, n_587);
  or g718 (n_675, wc3, n_579);
  not gc3 (wc3, n_580);
  or g719 (n_676, wc4, n_589);
  not gc4 (wc4, n_592);
  or g720 (n_677, wc5, n_594);
  not gc5 (wc5, n_597);
  or g721 (n_678, wc6, n_584);
  not gc6 (wc6, n_585);
  or g722 (n_679, wc7, n_599);
  not gc7 (wc7, n_602);
  or g723 (n_680, wc8, n_604);
  not gc8 (wc8, n_607);
  or g724 (n_681, wc9, n_589);
  not gc9 (wc9, n_590);
  or g725 (n_682, wc10, n_609);
  not gc10 (wc10, n_612);
  or g726 (n_683, wc11, n_614);
  not gc11 (wc11, n_617);
  or g727 (n_684, wc12, n_619);
  not gc12 (wc12, n_622);
  or g728 (n_685, wc13, n_624);
  not gc13 (wc13, n_627);
  or g729 (n_686, wc14, n_629);
  not gc14 (wc14, n_632);
  or g730 (n_687, wc15, n_634);
  not gc15 (wc15, n_637);
  or g731 (n_688, wc16, n_639);
  not gc16 (wc16, n_642);
  or g732 (n_689, wc17, n_644);
  not gc17 (wc17, n_647);
  or g733 (n_690, wc18, n_594);
  not gc18 (wc18, n_595);
  or g734 (n_691, wc19, n_599);
  not gc19 (wc19, n_600);
  or g735 (n_692, wc20, n_604);
  not gc20 (wc20, n_605);
  or g736 (n_693, wc21, n_609);
  not gc21 (wc21, n_610);
  or g737 (n_694, wc22, n_614);
  not gc22 (wc22, n_615);
  or g738 (n_695, wc23, n_619);
  not gc23 (wc23, n_620);
  or g739 (n_696, wc24, n_624);
  not gc24 (wc24, n_625);
  or g740 (n_697, wc25, n_629);
  not gc25 (wc25, n_630);
  or g741 (n_698, wc26, n_634);
  not gc26 (wc26, n_635);
  or g742 (n_699, wc27, n_639);
  not gc27 (wc27, n_640);
endmodule

module csa_tree_mul_25_40_group_52_GENERIC(in_0, in_1, out_0);
  input [15:0] in_0;
  input [7:0] in_1;
  output [16:0] out_0;
  wire [15:0] in_0;
  wire [7:0] in_1;
  wire [16:0] out_0;
  csa_tree_mul_25_40_group_52_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .out_0 (out_0));
endmodule

module mult_unsigned_GENERIC_REAL(A, B, Z);
// synthesis_equation "assign Z = $unsigned(A) * $unsigned(B);"
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_325;
  wire n_328, n_330, n_333, n_335, n_336, n_338, n_340, n_341;
  wire n_343, n_345, n_346, n_348, n_350, n_351, n_353, n_355;
  wire n_356, n_358, n_360, n_361, n_363, n_365, n_366, n_368;
  wire n_370, n_371, n_373, n_375, n_376, n_378, n_380, n_381;
  wire n_383, n_385, n_386, n_388, n_390, n_391, n_393, n_417;
  wire n_419, n_420, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445;
  and g1 (Z[0], A[0], B[0]);
  and g2 (n_46, A[1], B[0]);
  and g3 (n_63, A[2], B[0]);
  and g4 (n_67, A[3], B[0]);
  and g5 (n_72, A[4], B[0]);
  and g6 (n_80, A[5], B[0]);
  and g7 (n_90, A[6], B[0]);
  and g8 (n_103, A[7], B[0]);
  and g9 (n_61, A[0], B[1]);
  and g10 (n_45, A[1], B[1]);
  and g11 (n_68, A[2], B[1]);
  and g12 (n_73, A[3], B[1]);
  and g13 (n_64, A[4], B[1]);
  and g14 (n_91, A[5], B[1]);
  and g15 (n_104, A[6], B[1]);
  and g16 (n_120, A[7], B[1]);
  and g17 (n_66, A[0], B[2]);
  and g18 (n_70, A[1], B[2]);
  and g19 (n_76, A[2], B[2]);
  and g20 (n_83, A[3], B[2]);
  and g21 (n_94, A[4], B[2]);
  and g22 (n_108, A[5], B[2]);
  and g23 (n_121, A[6], B[2]);
  and g24 (n_137, A[7], B[2]);
  and g25 (n_69, A[0], B[3]);
  and g26 (n_74, A[1], B[3]);
  and g27 (n_81, A[2], B[3]);
  and g28 (n_92, A[3], B[3]);
  and g29 (n_105, A[4], B[3]);
  and g30 (n_124, A[5], B[3]);
  and g31 (n_138, A[6], B[3]);
  and g32 (n_152, A[7], B[3]);
  and g33 (n_75, A[0], B[4]);
  and g34 (n_82, A[1], B[4]);
  and g35 (n_93, A[2], B[4]);
  and g36 (n_107, A[3], B[4]);
  and g37 (n_122, A[4], B[4]);
  and g38 (n_141, A[5], B[4]);
  and g39 (n_153, A[6], B[4]);
  and g40 (n_164, A[7], B[4]);
  and g41 (n_84, A[0], B[5]);
  and g42 (n_65, A[1], B[5]);
  and g43 (n_109, A[2], B[5]);
  and g44 (n_123, A[3], B[5]);
  and g45 (n_139, A[4], B[5]);
  and g46 (n_156, A[5], B[5]);
  and g47 (n_165, A[6], B[5]);
  and g48 (n_173, A[7], B[5]);
  and g49 (n_95, A[0], B[6]);
  and g50 (n_110, A[1], B[6]);
  and g51 (n_125, A[2], B[6]);
  and g52 (n_140, A[3], B[6]);
  and g53 (n_154, A[4], B[6]);
  and g54 (n_167, A[5], B[6]);
  and g55 (n_174, A[6], B[6]);
  and g56 (n_179, A[7], B[6]);
  and g57 (n_106, A[0], B[7]);
  and g58 (n_126, A[1], B[7]);
  and g59 (n_142, A[2], B[7]);
  and g60 (n_155, A[3], B[7]);
  and g61 (n_166, A[4], B[7]);
  and g62 (n_175, A[5], B[7]);
  and g63 (n_180, A[6], B[7]);
  and g64 (n_33, A[7], B[7]);
  xor g107 (n_60, n_63, n_66);
  and g108 (n_44, n_63, n_66);
  xor g109 (n_71, n_67, n_68);
  and g110 (n_78, n_67, n_68);
  xor g111 (n_182, n_69, n_70);
  xor g112 (n_59, n_182, n_71);
  nand g113 (n_183, n_69, n_70);
  nand g114 (n_184, n_71, n_70);
  nand g115 (n_185, n_69, n_71);
  nand g116 (n_43, n_183, n_184, n_185);
  xor g117 (n_77, n_72, n_73);
  and g118 (n_86, n_72, n_73);
  xor g119 (n_186, n_74, n_75);
  xor g120 (n_79, n_186, n_76);
  nand g121 (n_187, n_74, n_75);
  nand g122 (n_188, n_76, n_75);
  nand g123 (n_189, n_74, n_76);
  nand g124 (n_87, n_187, n_188, n_189);
  xor g125 (n_190, n_77, n_78);
  xor g126 (n_58, n_190, n_79);
  nand g127 (n_191, n_77, n_78);
  nand g128 (n_192, n_79, n_78);
  nand g129 (n_193, n_77, n_79);
  nand g130 (n_42, n_191, n_192, n_193);
  xor g131 (n_85, n_80, n_64);
  and g132 (n_96, n_80, n_64);
  xor g133 (n_194, n_81, n_82);
  xor g134 (n_88, n_194, n_83);
  nand g135 (n_195, n_81, n_82);
  nand g136 (n_196, n_83, n_82);
  nand g137 (n_197, n_81, n_83);
  nand g138 (n_98, n_195, n_196, n_197);
  xor g139 (n_198, n_84, n_85);
  xor g140 (n_89, n_198, n_86);
  nand g141 (n_199, n_84, n_85);
  nand g142 (n_200, n_86, n_85);
  nand g143 (n_201, n_84, n_86);
  nand g144 (n_100, n_199, n_200, n_201);
  xor g145 (n_202, n_87, n_88);
  xor g146 (n_57, n_202, n_89);
  nand g147 (n_203, n_87, n_88);
  nand g148 (n_204, n_89, n_88);
  nand g149 (n_205, n_87, n_89);
  nand g150 (n_41, n_203, n_204, n_205);
  xor g151 (n_97, n_90, n_91);
  and g152 (n_111, n_90, n_91);
  xor g153 (n_206, n_92, n_93);
  xor g154 (n_99, n_206, n_94);
  nand g155 (n_207, n_92, n_93);
  nand g156 (n_208, n_94, n_93);
  nand g157 (n_209, n_92, n_94);
  nand g158 (n_113, n_207, n_208, n_209);
  xor g159 (n_210, n_65, n_95);
  xor g160 (n_101, n_210, n_96);
  nand g161 (n_211, n_65, n_95);
  nand g162 (n_212, n_96, n_95);
  nand g163 (n_213, n_65, n_96);
  nand g164 (n_116, n_211, n_212, n_213);
  xor g165 (n_214, n_97, n_98);
  xor g166 (n_102, n_214, n_99);
  nand g167 (n_215, n_97, n_98);
  nand g168 (n_216, n_99, n_98);
  nand g169 (n_217, n_97, n_99);
  nand g170 (n_118, n_215, n_216, n_217);
  xor g171 (n_218, n_100, n_101);
  xor g172 (n_56, n_218, n_102);
  nand g173 (n_219, n_100, n_101);
  nand g174 (n_220, n_102, n_101);
  nand g175 (n_221, n_100, n_102);
  nand g176 (n_40, n_219, n_220, n_221);
  xor g177 (n_112, n_103, n_104);
  and g178 (n_128, n_103, n_104);
  xor g179 (n_222, n_105, n_106);
  xor g180 (n_115, n_222, n_107);
  nand g181 (n_223, n_105, n_106);
  nand g182 (n_224, n_107, n_106);
  nand g183 (n_225, n_105, n_107);
  nand g184 (n_129, n_223, n_224, n_225);
  xor g185 (n_226, n_108, n_109);
  xor g186 (n_114, n_226, n_110);
  nand g187 (n_227, n_108, n_109);
  nand g188 (n_228, n_110, n_109);
  nand g189 (n_229, n_108, n_110);
  nand g190 (n_130, n_227, n_228, n_229);
  xor g191 (n_230, n_111, n_112);
  xor g192 (n_117, n_230, n_113);
  nand g193 (n_231, n_111, n_112);
  nand g194 (n_232, n_113, n_112);
  nand g195 (n_233, n_111, n_113);
  nand g196 (n_133, n_231, n_232, n_233);
  xor g197 (n_234, n_114, n_115);
  xor g198 (n_119, n_234, n_116);
  nand g199 (n_235, n_114, n_115);
  nand g200 (n_236, n_116, n_115);
  nand g201 (n_237, n_114, n_116);
  nand g202 (n_135, n_235, n_236, n_237);
  xor g203 (n_238, n_117, n_118);
  xor g204 (n_55, n_238, n_119);
  nand g205 (n_239, n_117, n_118);
  nand g206 (n_240, n_119, n_118);
  nand g207 (n_241, n_117, n_119);
  nand g208 (n_39, n_239, n_240, n_241);
  xor g209 (n_127, n_120, n_121);
  and g210 (n_143, n_120, n_121);
  xor g211 (n_242, n_122, n_123);
  xor g212 (n_131, n_242, n_124);
  nand g213 (n_243, n_122, n_123);
  nand g214 (n_244, n_124, n_123);
  nand g215 (n_245, n_122, n_124);
  nand g216 (n_144, n_243, n_244, n_245);
  xor g217 (n_246, n_125, n_126);
  xor g218 (n_132, n_246, n_127);
  nand g219 (n_247, n_125, n_126);
  nand g220 (n_248, n_127, n_126);
  nand g221 (n_249, n_125, n_127);
  nand g222 (n_147, n_247, n_248, n_249);
  xor g223 (n_250, n_128, n_129);
  xor g224 (n_134, n_250, n_130);
  nand g225 (n_251, n_128, n_129);
  nand g226 (n_252, n_130, n_129);
  nand g227 (n_253, n_128, n_130);
  nand g228 (n_148, n_251, n_252, n_253);
  xor g229 (n_254, n_131, n_132);
  xor g230 (n_136, n_254, n_133);
  nand g231 (n_255, n_131, n_132);
  nand g232 (n_256, n_133, n_132);
  nand g233 (n_257, n_131, n_133);
  nand g234 (n_151, n_255, n_256, n_257);
  xor g235 (n_258, n_134, n_135);
  xor g236 (n_54, n_258, n_136);
  nand g237 (n_259, n_134, n_135);
  nand g238 (n_260, n_136, n_135);
  nand g239 (n_261, n_134, n_136);
  nand g240 (n_38, n_259, n_260, n_261);
  xor g241 (n_262, n_137, n_138);
  xor g242 (n_146, n_262, n_139);
  nand g243 (n_263, n_137, n_138);
  nand g244 (n_264, n_139, n_138);
  nand g245 (n_265, n_137, n_139);
  nand g246 (n_158, n_263, n_264, n_265);
  xor g247 (n_266, n_140, n_141);
  xor g248 (n_145, n_266, n_142);
  nand g249 (n_267, n_140, n_141);
  nand g250 (n_268, n_142, n_141);
  nand g251 (n_269, n_140, n_142);
  nand g252 (n_157, n_267, n_268, n_269);
  xor g253 (n_270, n_143, n_144);
  xor g254 (n_149, n_270, n_145);
  nand g255 (n_271, n_143, n_144);
  nand g256 (n_272, n_145, n_144);
  nand g257 (n_273, n_143, n_145);
  nand g258 (n_161, n_271, n_272, n_273);
  xor g259 (n_274, n_146, n_147);
  xor g260 (n_150, n_274, n_148);
  nand g261 (n_275, n_146, n_147);
  nand g262 (n_276, n_148, n_147);
  nand g263 (n_277, n_146, n_148);
  nand g264 (n_163, n_275, n_276, n_277);
  xor g265 (n_278, n_149, n_150);
  xor g266 (n_53, n_278, n_151);
  nand g267 (n_279, n_149, n_150);
  nand g268 (n_280, n_151, n_150);
  nand g269 (n_281, n_149, n_151);
  nand g270 (n_37, n_279, n_280, n_281);
  xor g271 (n_282, n_152, n_153);
  xor g272 (n_159, n_282, n_154);
  nand g273 (n_283, n_152, n_153);
  nand g274 (n_284, n_154, n_153);
  nand g275 (n_285, n_152, n_154);
  nand g276 (n_168, n_283, n_284, n_285);
  xor g277 (n_286, n_155, n_156);
  xor g278 (n_160, n_286, n_157);
  nand g279 (n_287, n_155, n_156);
  nand g280 (n_288, n_157, n_156);
  nand g281 (n_289, n_155, n_157);
  nand g282 (n_170, n_287, n_288, n_289);
  xor g283 (n_290, n_158, n_159);
  xor g284 (n_162, n_290, n_160);
  nand g285 (n_291, n_158, n_159);
  nand g286 (n_292, n_160, n_159);
  nand g287 (n_293, n_158, n_160);
  nand g288 (n_172, n_291, n_292, n_293);
  xor g289 (n_294, n_161, n_162);
  xor g290 (n_52, n_294, n_163);
  nand g291 (n_295, n_161, n_162);
  nand g292 (n_296, n_163, n_162);
  nand g293 (n_297, n_161, n_163);
  nand g294 (n_36, n_295, n_296, n_297);
  xor g295 (n_298, n_164, n_165);
  xor g296 (n_169, n_298, n_166);
  nand g297 (n_299, n_164, n_165);
  nand g298 (n_300, n_166, n_165);
  nand g299 (n_301, n_164, n_166);
  nand g300 (n_176, n_299, n_300, n_301);
  xor g301 (n_302, n_167, n_168);
  xor g302 (n_171, n_302, n_169);
  nand g303 (n_303, n_167, n_168);
  nand g304 (n_304, n_169, n_168);
  nand g305 (n_305, n_167, n_169);
  nand g306 (n_178, n_303, n_304, n_305);
  xor g307 (n_306, n_170, n_171);
  xor g308 (n_51, n_306, n_172);
  nand g309 (n_307, n_170, n_171);
  nand g310 (n_308, n_172, n_171);
  nand g311 (n_309, n_170, n_172);
  nand g312 (n_50, n_307, n_308, n_309);
  xor g313 (n_310, n_173, n_174);
  xor g314 (n_177, n_310, n_175);
  nand g315 (n_311, n_173, n_174);
  nand g316 (n_312, n_175, n_174);
  nand g317 (n_313, n_173, n_175);
  nand g318 (n_181, n_311, n_312, n_313);
  xor g319 (n_314, n_176, n_177);
  xor g320 (n_35, n_314, n_178);
  nand g321 (n_315, n_176, n_177);
  nand g322 (n_316, n_178, n_177);
  nand g323 (n_317, n_176, n_178);
  nand g324 (n_49, n_315, n_316, n_317);
  xor g325 (n_318, n_179, n_180);
  xor g326 (n_34, n_318, n_181);
  nand g327 (n_319, n_179, n_180);
  nand g328 (n_320, n_181, n_180);
  nand g329 (n_321, n_179, n_181);
  nand g330 (n_48, n_319, n_320, n_321);
  nor g336 (n_325, n_46, n_61);
  nand g337 (n_328, n_46, n_61);
  nor g338 (n_330, n_45, n_60);
  nand g339 (n_333, n_45, n_60);
  nor g340 (n_335, n_44, n_59);
  nand g341 (n_338, n_44, n_59);
  nor g342 (n_340, n_43, n_58);
  nand g343 (n_343, n_43, n_58);
  nor g344 (n_345, n_42, n_57);
  nand g345 (n_348, n_42, n_57);
  nor g346 (n_350, n_41, n_56);
  nand g347 (n_353, n_41, n_56);
  nor g348 (n_355, n_40, n_55);
  nand g349 (n_358, n_40, n_55);
  nor g350 (n_360, n_39, n_54);
  nand g351 (n_363, n_39, n_54);
  nor g352 (n_365, n_38, n_53);
  nand g353 (n_368, n_38, n_53);
  nor g354 (n_370, n_37, n_52);
  nand g355 (n_373, n_37, n_52);
  nor g356 (n_375, n_36, n_51);
  nand g357 (n_378, n_36, n_51);
  nor g358 (n_380, n_35, n_50);
  nand g359 (n_383, n_35, n_50);
  nor g360 (n_385, n_34, n_49);
  nand g361 (n_388, n_34, n_49);
  nor g362 (n_390, n_33, n_48);
  nand g363 (n_393, n_33, n_48);
  nand g371 (n_336, n_333, n_420);
  nand g374 (n_341, n_338, n_424);
  nand g377 (n_346, n_343, n_428);
  nand g380 (n_351, n_348, n_434);
  nand g383 (n_356, n_353, n_437);
  nand g386 (n_361, n_358, n_438);
  nand g389 (n_366, n_363, n_439);
  nand g392 (n_371, n_368, n_440);
  nand g65 (n_376, n_373, n_441);
  nand g68 (n_381, n_378, n_442);
  nand g71 (n_386, n_383, n_443);
  nand g74 (n_391, n_388, n_444);
  nand g77 (Z[15], n_393, n_445);
  xnor g86 (Z[3], n_336, n_422);
  xnor g88 (Z[4], n_341, n_423);
  xnor g90 (Z[5], n_346, n_425);
  xnor g92 (Z[6], n_351, n_427);
  xnor g94 (Z[7], n_356, n_429);
  xnor g96 (Z[8], n_361, n_431);
  xnor g98 (Z[9], n_366, n_432);
  xnor g100 (Z[10], n_371, n_435);
  xnor g102 (Z[11], n_376, n_436);
  xnor g104 (Z[12], n_381, n_433);
  xnor g106 (Z[13], n_386, n_430);
  xnor g396 (Z[14], n_391, n_426);
  or g400 (n_417, wc, n_325);
  not gc (wc, n_328);
  not g402 (Z[1], n_417);
  or g403 (n_419, wc0, n_330);
  not gc0 (wc0, n_333);
  or g404 (n_420, n_328, n_330);
  xor g405 (Z[2], n_328, n_419);
  or g406 (n_422, wc1, n_335);
  not gc1 (wc1, n_338);
  or g407 (n_423, wc2, n_340);
  not gc2 (wc2, n_343);
  or g408 (n_424, wc3, n_335);
  not gc3 (wc3, n_336);
  or g409 (n_425, wc4, n_345);
  not gc4 (wc4, n_348);
  or g410 (n_426, wc5, n_390);
  not gc5 (wc5, n_393);
  or g411 (n_427, wc6, n_350);
  not gc6 (wc6, n_353);
  or g412 (n_428, wc7, n_340);
  not gc7 (wc7, n_341);
  or g413 (n_429, wc8, n_355);
  not gc8 (wc8, n_358);
  or g414 (n_430, wc9, n_385);
  not gc9 (wc9, n_388);
  or g415 (n_431, wc10, n_360);
  not gc10 (wc10, n_363);
  or g416 (n_432, wc11, n_365);
  not gc11 (wc11, n_368);
  or g417 (n_433, wc12, n_380);
  not gc12 (wc12, n_383);
  or g418 (n_434, wc13, n_345);
  not gc13 (wc13, n_346);
  or g419 (n_435, wc14, n_370);
  not gc14 (wc14, n_373);
  or g420 (n_436, wc15, n_375);
  not gc15 (wc15, n_378);
  or g421 (n_437, wc16, n_350);
  not gc16 (wc16, n_351);
  or g422 (n_438, wc17, n_355);
  not gc17 (wc17, n_356);
  or g423 (n_439, wc18, n_360);
  not gc18 (wc18, n_361);
  or g424 (n_440, wc19, n_365);
  not gc19 (wc19, n_366);
  or g425 (n_441, wc20, n_370);
  not gc20 (wc20, n_371);
  or g426 (n_442, wc21, n_375);
  not gc21 (wc21, n_376);
  or g427 (n_443, wc22, n_380);
  not gc22 (wc22, n_381);
  or g428 (n_444, wc23, n_385);
  not gc23 (wc23, n_386);
  or g429 (n_445, wc24, n_390);
  not gc24 (wc24, n_391);
endmodule

module mult_unsigned_GENERIC(A, B, Z);
  input [7:0] A, B;
  output [15:0] Z;
  wire [7:0] A, B;
  wire [15:0] Z;
  mult_unsigned_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

