###############################################################################
#TSMC Library/IP Product
#Filename: tcbn65gplus_8lmT2.lef
#Technology: CLN65GPLUS
#Product Type: Standard Cell
#Product Name: tcbn65gplus
#Version: 121a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

# DESIGN RULE DOCUMENT: T-N65-CL-DR-001 V1.2
# SPICE MODEL DOCUMENT: T-N65-CL-SP-031 V1.0
# Resistor & Capacitor are referenced from spice model interconnect table
# The index is "width=minWidth", "Space=Pitch"
VERSION	5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
    CAPACITANCE PICOFARADS 10 ;
    CURRENT MILLIAMPS 10000 ;
    VOLTAGE VOLTS 1000 ;
    FREQUENCY MEGAHERTZ 10 ;
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER PO
    TYPE MASTERSLICE ;
END PO

LAYER CO
    TYPE CUT ;
END CO

PROPERTYDEFINITIONS 
    LAYER LEF57_SPACING STRING ;
END PROPERTYDEFINITIONS 

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    OFFSET 0.000 ;
    HEIGHT 0.5900 ;
    THICKNESS 0.1800 ;
    MINSTEP 0.090 ; 
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.09 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.42    1.50    4.50
    WIDTH    0.00         0.09    0.09    0.09    0.09    0.09
    WIDTH    0.20         0.09    0.11    0.11    0.11    0.11
    WIDTH    0.42         0.09    0.11    0.16    0.16    0.16
    WIDTH    1.50         0.09    0.11    0.16    0.50    0.50
    WIDTH    4.50         0.09    0.11    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.11 ENDOFLINE 0.11 WITHIN 0.035 PARALLELEDGE 0.11 WITHIN 0.11 ;" ;
    AREA 0.042 ;
    MINENCLOSEDAREA 0.20 ;

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;

    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.801 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.001 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.001 ;

    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

    ACCURRENTDENSITY 	AVERAGE
        FREQUENCY 	500 ;
        WIDTH     	0.090 	1.000 ;
        TABLEENTRIES	1.241	1.485 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH		0.090	0.180	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	14.936	13.727	11.656	10.736	9.829	9.681 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.090 1.0 12 ;
        TABLEENTRIES	41.861 50.097 50.844 ;
    RESISTANCE RPERSQ 0.1600000000 ;
    CAPACITANCE CPERSQDIST 0.0001711111 ;
    EDGECAPACITANCE 0.0000883000 ;
END M1

LAYER VIA1
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA1

LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    OFFSET 0.100 ;
    HEIGHT 0.9450 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;

    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.801 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.001 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.001 ;

    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	9.324	8.384	7.101	6.451	5.803	5.696 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;
                		
    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000780000 ;
END M2

LAYER VIA2
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA2

LAYER M3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    OFFSET 0.000 ;
    HEIGHT 1.3400 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;

    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.801 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.001 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.001 ;

    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.965	7.789	6.191	5.347	4.453	4.299 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;
              		
    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000779000 ;
END M3

LAYER VIA3
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA3

LAYER M4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    OFFSET 0.100 ;
    HEIGHT 1.7350 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.801 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.001 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.824	7.548	5.805	4.857	3.811	3.623 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;

    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000778000 ;
END M4

LAYER VIA4
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA4

LAYER M5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    OFFSET 0.000 ;
    HEIGHT 2.1300 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.801 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.001 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.752	7.421	5.592	4.578	3.423	3.208 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;

    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000778000 ;
END M5

LAYER VIA5
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA5

LAYER M6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    OFFSET 0.100 ;
    HEIGHT 2.5250 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 0.300 FROMBELOW ;
    MINIMUMCUT 4 WIDTH 0.700 FROMBELOW ;
    MINIMUMCUT 2 WIDTH 0.300 FROMBELOW LENGTH 0.300 WITHIN 0.801 ;
    MINIMUMCUT 2 WIDTH 2.000 FROMBELOW LENGTH 2.000 WITHIN 2.001 ;
    MINIMUMCUT 2 WIDTH 3.000 FROMBELOW LENGTH 10.000 WITHIN 5.001 ;
    MINIMUMCUT 2 WIDTH 1.800 FROMABOVE ;
    MINIMUMCUT 2 WIDTH 3.000 FROMABOVE LENGTH 10.0 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100   1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.701	7.336	5.453	4.394	3.158	2.921 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;

    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000778000 ;
END M6

LAYER VIA6
    TYPE CUT ;
    SPACING 0.340 ;
    SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	23.742 ;
END VIA6

LAYER M7
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.800 ;
    OFFSET 0.000 ;
    HEIGHT 3.3400 ;
    THICKNESS 0.9000 ;
    MINSTEP 0.400 ;
    FILLACTIVESPACING 0.600 ;
    WIDTH 0.400 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    1.50    4.50
    WIDTH    0.00         0.40    0.40    0.40
    WIDTH    1.50         0.40    0.50    0.50
    WIDTH    4.50         0.40    0.50    1.50 ;
    AREA 0.565 ;
    MINENCLOSEDAREA 0.565 ;   

    MINIMUMDENSITY 20 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 80 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;

    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 1.800 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.0 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.400	1.000 ;
        TABLEENTRIES 	7.691	7.934 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.400	0.600	0.800	1.000	5.000	12.000 ;
        TABLEENTRIES	11.490	9.972	9.037	8.396	5.667	5.116 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.400 1.0 12 ;
        TABLEENTRIES	84.641 87.314 88.947 ;
  
    RESISTANCE RPERSQ 0.0220000000 ;
    CAPACITANCE CPERSQDIST 0.0000632500 ;
    EDGECAPACITANCE 0.0000915000 ;
END M7

LAYER VIA7
    TYPE CUT ;
    SPACING 0.340 ;
    SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	23.742 ;
END VIA7

LAYER M8
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.800 ;
    OFFSET 0.100 ;
    HEIGHT 4.8350 ;
    THICKNESS 0.9000 ;
    MINSTEP 0.400 ;
    FILLACTIVESPACING 0.600 ;
    WIDTH 0.400 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    1.50    4.50
    WIDTH    0.00         0.40    0.40    0.40
    WIDTH    1.50         0.40    0.50    0.50
    WIDTH    4.50         0.40    0.50    1.50 ;
    AREA 0.565 ;
    MINENCLOSEDAREA 0.565 ;   

    MINIMUMDENSITY 20 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 80 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;

    MINIMUMDENSITY 1 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 1.800 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.0 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 50480 ) ( 0.5 54000 ) ( 1 58000 ) ( 1.5 62000 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.400	1.000 ;
        TABLEENTRIES 	7.691	7.934 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.400	0.600	0.800	1.000	5.000	12.000 ;
        TABLEENTRIES	11.373	9.827	8.870	8.213	5.372	4.783 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.400 1.0 12 ;
        TABLEENTRIES	84.641 87.314 88.947 ;

    RESISTANCE RPERSQ 0.0220000000 ;
    CAPACITANCE CPERSQDIST 0.0000632500 ;
    EDGECAPACITANCE 0.0000956000 ;
END M8

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA12_1cut

VIA VIA12_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA12_1cut_H
                 
VIA VIA12_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA12_1cut_V

VIA VIA12_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA12_1cut_FAT_C
             
VIA VIA12_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA12_1cut_FAT_H

VIA VIA12_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA12_1cut_FAT_V

VIA VIA12_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA12_1cut_FAT
                 
VIA VIA12_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA12_2cut_E

VIA VIA12_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M2 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA12_2cut_W

VIA VIA12_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA12_2cut_N

VIA VIA12_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M2 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA12_2cut_S

VIA VIA12_2cut_HN DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.050 -0.090  0.050  0.330 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.190  0.050  0.290 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.330 ;
END VIA12_2cut_HN

VIA VIA12_2cut_HS DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.050 -0.330  0.050  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.290  0.050 -0.190 ;
    LAYER M2 ;
        RECT -0.050 -0.330  0.050  0.090 ;
END VIA12_2cut_HS

VIA VIA12_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M1 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA1 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M2 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA12_4cut

VIA VIA23_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1cut

VIA VIA23_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA23_1cut_V
                 
VIA VIA23_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1cut_H

VIA VIA23_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA23_1cut_FAT_C
             
VIA VIA23_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA23_1cut_FAT_V

VIA VIA23_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA23_1cut_FAT_H

VIA VIA23_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA23_1cut_FAT
                 
VIA VIA23_1stack_N DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.430 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1stack_N

VIA VIA23_1stack_S DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.430  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1stack_S

VIA VIA23_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.250  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.290  0.050 ;
END VIA23_2cut_E

VIA VIA23_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.250 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M3 ;
        RECT -0.290 -0.050  0.090  0.050 ;
END VIA23_2cut_W

VIA VIA23_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.290 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.250 ;
END VIA23_2cut_N

VIA VIA23_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.050 -0.290  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M3 ;
        RECT -0.090 -0.250  0.090  0.050 ;
END VIA23_2cut_S

VIA VIA23_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M2 ;
        RECT -0.150 -0.190  0.150  0.190 ;
    LAYER VIA2 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M3 ;
        RECT -0.190 -0.150  0.190  0.150 ;
END VIA23_4cut

VIA VIA34_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1cut

VIA VIA34_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA34_1cut_H
                 
VIA VIA34_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1cut_V

VIA VIA34_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA34_1cut_FAT_C
             
VIA VIA34_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA34_1cut_FAT_H

VIA VIA34_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA34_1cut_FAT_V

VIA VIA34_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA34_1cut_FAT
                 
VIA VIA34_1stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.430  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1stack_E

VIA VIA34_1stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.430 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1stack_W

VIA VIA34_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA34_2cut_E

VIA VIA34_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M4 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA34_2cut_W

VIA VIA34_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA34_2cut_N

VIA VIA34_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M4 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA34_2cut_S

VIA VIA34_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M3 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA3 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M4 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA34_4cut

VIA VIA45_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1cut

VIA VIA45_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA45_1cut_V
                 
VIA VIA45_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1cut_H

VIA VIA45_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA45_1cut_FAT_C
             
VIA VIA45_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA45_1cut_FAT_V

VIA VIA45_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA45_1cut_FAT_H

VIA VIA45_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA45_1cut_FAT
                 
VIA VIA45_1stack_N DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.430 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1stack_N

VIA VIA45_1stack_S DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.430  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1stack_S

VIA VIA45_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.250  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.290  0.050 ;
END VIA45_2cut_E

VIA VIA45_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.250 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M5 ;
        RECT -0.290 -0.050  0.090  0.050 ;
END VIA45_2cut_W

VIA VIA45_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.290 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.250 ;
END VIA45_2cut_N

VIA VIA45_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.050 -0.290  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M5 ;
        RECT -0.090 -0.250  0.090  0.050 ;
END VIA45_2cut_S

VIA VIA45_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M4 ;
        RECT -0.150 -0.190  0.150  0.190 ;
    LAYER VIA4 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M5 ;
        RECT -0.190 -0.150  0.190  0.150 ;
END VIA45_4cut

VIA VIA56_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1cut

VIA VIA56_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA56_1cut_H
                 
VIA VIA56_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1cut_V

VIA VIA56_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA56_1cut_FAT_C
             
VIA VIA56_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA56_1cut_FAT_H

VIA VIA56_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA56_1cut_FAT_V

VIA VIA56_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA56_1cut_FAT
                 
VIA VIA56_1stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.430  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1stack_E

VIA VIA56_1stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.430 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1stack_W

VIA VIA56_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA56_2cut_E

VIA VIA56_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M6 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA56_2cut_W

VIA VIA56_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA56_2cut_N

VIA VIA56_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M6 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA56_2cut_S

VIA VIA56_2stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.430  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA56_2stack_E
 
VIA VIA56_2stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.430 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M6 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA56_2stack_W

VIA VIA56_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M5 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA5 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M6 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA56_4cut

VIA VIA67_1cut DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut
 
VIA VIA67_1cut_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA67_1cut_V
 
VIA VIA67_1cut_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut_H
 
VIA VIA67_1cut_FAT_C DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.26  0.200  0.26 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
END VIA67_1cut_FAT_C
 
VIA VIA67_1cut_FAT_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.26  0.200  0.26 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA67_1cut_FAT_V
 
VIA VIA67_1cut_FAT_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
END VIA67_1cut_FAT_H
 
VIA VIA67_1cut_FAT DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.260 -0.260  0.260  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.260  0.260  0.260 ;
END VIA67_1cut_FAT
 
VIA VIA67_2cut_E DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.900  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT  0.520 -0.180  0.880  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.960  0.200 ;
END VIA67_2cut_E
 
VIA VIA67_2cut_W DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.900 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180 -0.520  0.180 ;
    LAYER M7 ;
        RECT -0.960 -0.200  0.260  0.200 ;
END VIA67_2cut_W
 
VIA VIA67_2cut_N DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.960 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180  0.520  0.180  0.880 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.900 ;
END VIA67_2cut_N
 
VIA VIA67_2cut_S DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.200 -0.960  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 -0.880  0.180 -0.520 ;
    LAYER M7 ;
        RECT -0.260 -0.900  0.260  0.200 ;
END VIA67_2cut_S
 
VIA VIA67_4cut DEFAULT
    RESISTANCE 0.0550000000 ;
    LAYER M6 ;
        RECT -0.650 -0.710  0.650  0.710 ;
    LAYER VIA6 ;
        RECT -0.630 -0.630 -0.270 -0.270 ;
        RECT -0.630  0.270 -0.270  0.630 ;
        RECT  0.270  0.270  0.630  0.630 ;
        RECT  0.270 -0.630  0.630 -0.270 ;
    LAYER M7 ;
        RECT -0.710 -0.650  0.710  0.650 ;
END VIA67_4cut

VIA VIA78_1cut DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut
 
VIA VIA78_1cut_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA78_1cut_H
 
VIA VIA78_1cut_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut_V
 
VIA VIA78_1cut_FAT_C DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA78_1cut_FAT_C
 
VIA VIA78_1cut_FAT_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.26 -0.200  0.26  0.200 ;
END VIA78_1cut_FAT_H
 
VIA VIA78_1cut_FAT_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.200 -0.26  0.200  0.26 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA78_1cut_FAT_V
 
VIA VIA78_1cut_FAT DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.260  0.260  0.260 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.260 -0.260  0.260  0.260 ;
END VIA78_1cut_FAT

VIA VIA78_1stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  1.155  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1stack_E
 
VIA VIA78_1stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -1.155 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1stack_W
 
VIA VIA78_2cut_E DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.960  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT  0.520 -0.180  0.880  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.900  0.260 ;
END VIA78_2cut_E
 
VIA VIA78_2cut_W DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.960 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180 -0.520  0.180 ;
    LAYER M8 ;
        RECT -0.900 -0.260  0.200  0.260 ;
END VIA78_2cut_W
 
VIA VIA78_2cut_N DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.900 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180  0.520  0.180  0.880 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.960 ;
END VIA78_2cut_N
 
VIA VIA78_2cut_S DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.260 -0.900  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 -0.880  0.180 -0.520 ;
    LAYER M8 ;
        RECT -0.200 -0.960  0.200  0.260 ;
END VIA78_2cut_S
 
VIA VIA78_4cut DEFAULT
    RESISTANCE 0.0550000000 ;
    LAYER M7 ;
        RECT -0.710 -0.650  0.710  0.650 ;
    LAYER VIA7 ;
        RECT -0.630 -0.630 -0.270 -0.270 ;
        RECT -0.630  0.270 -0.270  0.630 ;
        RECT  0.270  0.270  0.630  0.630 ;
        RECT  0.270 -0.630  0.630 -0.270 ;
    LAYER M8 ;
        RECT -0.650 -0.710  0.650  0.710 ;
END VIA78_4cut
 
VIARULE VIAGEN12 GENERATE
    LAYER M1 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.09 TO 12.00 ;
    LAYER M2 ;
        ENCLOSURE 0.4E-01 0 ;
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA1 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ;
        SPACING 0.23 BY 0.23 ;    
END VIAGEN12        

VIARULE VIAGEN23 GENERATE
    LAYER M2 ;
        ENCLOSURE 0.4E-01 0 ;  
        WIDTH 0.10 TO 12.00 ;
    LAYER M3 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA2 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN23

VIARULE VIAGEN34 GENERATE
    LAYER M3 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M4 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA3 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN34

VIARULE VIAGEN45 GENERATE
    LAYER M4 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M5 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA4 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN45

VIARULE VIAGEN56 GENERATE
    LAYER M5 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M6 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA5 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN56

VIARULE VIAGEN67 GENERATE
    LAYER M6 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.10 TO 12.00 ;
    LAYER M7 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.40 TO 12.00 ;
    LAYER VIA6 ;
        RECT -0.18 -0.18 0.18 0.18 ; 
        SPACING 0.90 BY 0.90 ;    
END VIAGEN67

VIARULE VIAGEN78 GENERATE
    LAYER M7 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.40 TO 12.00 ;
    LAYER M8 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.40 TO 12.00 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ; 
        SPACING 0.90 BY 0.90 ;    
END VIAGEN78           

MAXVIASTACK 4 RANGE M1 M6 ;

VIARULE TURN1 GENERATE
    LAYER M1 ;
        DIRECTION HORIZONTAL ;
    LAYER M1 ;
        DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
    LAYER M2 ;
        DIRECTION HORIZONTAL ;
    LAYER M2 ;
        DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
    LAYER M3 ;
        DIRECTION HORIZONTAL ;
    LAYER M3 ;
        DIRECTION VERTICAL ;
END TURN3

VIARULE TURN4 GENERATE
    LAYER M4 ;
        DIRECTION HORIZONTAL ;
    LAYER M4 ;
        DIRECTION VERTICAL ;
END TURN4

VIARULE TURN5 GENERATE
    LAYER M5 ;
        DIRECTION HORIZONTAL ;
    LAYER M5 ;
        DIRECTION VERTICAL ;
END TURN5

VIARULE TURN6 GENERATE
    LAYER M6 ;
        DIRECTION HORIZONTAL ;
    LAYER M6 ;
        DIRECTION VERTICAL ;
END TURN6

VIARULE TURN7 GENERATE
    LAYER M7 ;
        DIRECTION HORIZONTAL ;
    LAYER M7 ;
        DIRECTION VERTICAL ;
END TURN7

VIARULE TURN8 GENERATE
    LAYER M8 ;
        DIRECTION HORIZONTAL ;
    LAYER M8 ;
        DIRECTION VERTICAL ;
END TURN8

SITE core
    SIZE 0.20 BY 1.80 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END core

SITE bcore
    SIZE 0.20 BY 3.60 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END bcore
 
SITE ccore
    SIZE 0.20 BY 5.40 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END ccore
 
SITE dcore
    SIZE 0.20 BY 7.20 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END dcore
 
SITE gacore
    SIZE 0.80 BY 1.80 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END gacore

MACRO AN2D0
    CLASS CORE ;
    FOREIGN AN2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.285 1.150 1.490 ;
        RECT  0.980 0.285 1.050 0.475 ;
        RECT  0.980 1.060 1.050 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.680 0.640 0.930 ;
        RECT  0.450 0.680 0.550 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 -0.165 1.200 0.165 ;
        RECT  0.670 -0.165 0.820 0.360 ;
        RECT  0.000 -0.165 0.670 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.635 1.200 1.965 ;
        RECT  0.690 1.440 0.800 1.965 ;
        RECT  0.225 1.635 0.690 1.965 ;
        RECT  0.105 1.240 0.225 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.870 0.750 0.930 0.940 ;
        RECT  0.760 0.470 0.870 1.330 ;
        RECT  0.485 0.470 0.760 0.570 ;
        RECT  0.340 1.230 0.760 1.330 ;
        RECT  0.375 0.320 0.485 0.570 ;
        RECT  0.090 0.320 0.375 0.450 ;
    END
END AN2D0

MACRO AN2D1
    CLASS CORE ;
    FOREIGN AN2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.285 1.150 1.490 ;
        RECT  0.980 0.285 1.050 0.475 ;
        RECT  0.980 1.060 1.050 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.680 0.640 0.930 ;
        RECT  0.450 0.680 0.550 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 -0.165 1.200 0.165 ;
        RECT  0.670 -0.165 0.820 0.360 ;
        RECT  0.000 -0.165 0.670 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.635 1.200 1.965 ;
        RECT  0.670 1.440 0.820 1.965 ;
        RECT  0.225 1.635 0.670 1.965 ;
        RECT  0.105 1.230 0.225 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.870 0.750 0.930 0.940 ;
        RECT  0.760 0.470 0.870 1.330 ;
        RECT  0.485 0.470 0.760 0.570 ;
        RECT  0.340 1.230 0.760 1.330 ;
        RECT  0.375 0.320 0.485 0.570 ;
        RECT  0.090 0.320 0.375 0.450 ;
    END
END AN2D1

MACRO AN2D2
    CLASS CORE ;
    FOREIGN AN2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.545 1.150 1.195 ;
        RECT  0.940 0.275 1.050 0.675 ;
        RECT  1.040 1.045 1.050 1.195 ;
        RECT  0.930 1.045 1.040 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.680 0.600 0.930 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.100 ;
        RECT  0.210 0.680 0.250 0.950 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 -0.165 1.400 0.165 ;
        RECT  1.195 -0.165 1.315 0.455 ;
        RECT  0.785 -0.165 1.195 0.165 ;
        RECT  0.635 -0.165 0.785 0.350 ;
        RECT  0.000 -0.165 0.635 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 1.635 1.400 1.965 ;
        RECT  1.195 1.335 1.315 1.965 ;
        RECT  0.225 1.635 1.195 1.965 ;
        RECT  0.225 1.390 0.820 1.490 ;
        RECT  0.105 1.210 0.225 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.820 0.775 0.930 0.945 ;
        RECT  0.720 0.460 0.820 1.300 ;
        RECT  0.080 0.460 0.720 0.570 ;
        RECT  0.340 1.210 0.720 1.300 ;
    END
END AN2D2

MACRO AN2D4
    CLASS CORE ;
    FOREIGN AN2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.435 2.100 0.615 ;
        RECT  1.850 1.110 2.100 1.290 ;
        RECT  1.550 0.435 1.850 1.290 ;
        RECT  1.390 0.435 1.550 0.615 ;
        RECT  1.390 1.110 1.550 1.290 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.975 0.665 1.090 0.940 ;
        RECT  0.760 0.665 0.975 0.765 ;
        RECT  0.650 0.500 0.760 0.765 ;
        RECT  0.360 0.500 0.650 0.590 ;
        RECT  0.270 0.500 0.360 0.780 ;
        RECT  0.190 0.680 0.270 0.780 ;
        RECT  0.050 0.680 0.190 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.900 0.750 1.100 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.165 2.400 0.165 ;
        RECT  2.210 -0.165 2.330 0.705 ;
        RECT  1.820 -0.165 2.210 0.165 ;
        RECT  1.630 -0.165 1.820 0.325 ;
        RECT  1.225 -0.165 1.630 0.165 ;
        RECT  1.075 -0.165 1.225 0.345 ;
        RECT  0.180 -0.165 1.075 0.165 ;
        RECT  0.060 -0.165 0.180 0.570 ;
        RECT  0.000 -0.165 0.060 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.635 2.400 1.965 ;
        RECT  2.210 1.095 2.330 1.965 ;
        RECT  1.170 1.635 2.210 1.965 ;
        RECT  1.170 1.390 1.830 1.490 ;
        RECT  1.030 1.390 1.170 1.965 ;
        RECT  0.550 1.390 1.030 1.490 ;
        RECT  0.190 1.635 1.030 1.965 ;
        RECT  0.070 1.230 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.950 0.435 2.100 0.615 ;
        RECT  1.950 1.110 2.100 1.290 ;
        RECT  1.390 0.435 1.450 0.615 ;
        RECT  1.390 1.110 1.450 1.290 ;
        RECT  1.290 0.730 1.405 0.940 ;
        RECT  1.190 0.455 1.290 1.300 ;
        RECT  0.950 0.455 1.190 0.555 ;
        RECT  0.300 1.210 1.190 1.300 ;
        RECT  0.850 0.310 0.950 0.555 ;
        RECT  0.525 0.310 0.850 0.410 ;
    END
END AN2D4

MACRO AN2D8
    CLASS CORE ;
    FOREIGN AN2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.310 3.505 0.690 ;
        RECT  2.850 1.110 3.505 1.490 ;
        RECT  2.550 0.310 2.850 1.490 ;
        RECT  1.840 0.310 2.550 0.690 ;
        RECT  1.840 1.110 2.550 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.570 1.550 0.955 ;
        RECT  0.750 0.570 1.435 0.660 ;
        RECT  0.650 0.570 0.750 0.900 ;
        RECT  0.450 0.700 0.650 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.750 1.165 1.120 ;
        RECT  0.190 1.020 1.035 1.120 ;
        RECT  0.050 0.700 0.190 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.735 -0.165 3.800 0.165 ;
        RECT  3.615 -0.165 3.735 0.690 ;
        RECT  0.730 -0.165 3.615 0.165 ;
        RECT  0.560 -0.165 0.730 0.300 ;
        RECT  0.000 -0.165 0.560 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.735 1.635 3.800 1.965 ;
        RECT  3.615 1.110 3.735 1.965 ;
        RECT  1.245 1.635 3.615 1.965 ;
        RECT  1.055 1.395 1.245 1.965 ;
        RECT  0.185 1.635 1.055 1.965 ;
        RECT  0.065 1.250 0.185 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.310 3.505 0.690 ;
        RECT  2.950 1.110 3.505 1.490 ;
        RECT  1.840 0.310 2.450 0.690 ;
        RECT  1.840 1.110 2.450 1.490 ;
        RECT  1.750 0.800 2.410 0.900 ;
        RECT  1.660 0.390 1.750 1.305 ;
        RECT  0.050 0.390 1.660 0.480 ;
        RECT  0.295 1.215 1.660 1.305 ;
    END
END AN2D8

MACRO AN2XD1
    CLASS CORE ;
    FOREIGN AN2XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.285 1.150 1.490 ;
        RECT  0.980 0.285 1.050 0.475 ;
        RECT  0.980 1.060 1.050 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.680 0.640 0.930 ;
        RECT  0.450 0.680 0.550 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 -0.165 1.200 0.165 ;
        RECT  0.670 -0.165 0.820 0.360 ;
        RECT  0.000 -0.165 0.670 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.635 1.200 1.965 ;
        RECT  0.670 1.440 0.820 1.965 ;
        RECT  0.225 1.635 0.670 1.965 ;
        RECT  0.105 1.230 0.225 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.870 0.750 0.930 0.940 ;
        RECT  0.760 0.460 0.870 1.330 ;
        RECT  0.080 0.460 0.760 0.570 ;
        RECT  0.340 1.230 0.760 1.330 ;
    END
END AN2XD1

MACRO AN3D0
    CLASS CORE ;
    FOREIGN AN3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.275 1.350 1.330 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.680 0.950 1.120 ;
        RECT  0.780 0.680 0.850 0.930 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.680 0.610 0.910 ;
        RECT  0.450 0.680 0.550 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.165 1.400 0.165 ;
        RECT  0.880 -0.165 1.070 0.300 ;
        RECT  0.000 -0.165 0.880 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.635 1.400 1.965 ;
        RECT  0.880 1.460 1.070 1.965 ;
        RECT  0.585 1.635 0.880 1.965 ;
        RECT  0.395 1.460 0.585 1.965 ;
        RECT  0.000 1.635 0.395 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.045 0.410 1.135 1.350 ;
        RECT  0.100 0.410 1.045 0.520 ;
        RECT  0.760 1.230 1.045 1.350 ;
        RECT  0.650 1.075 0.760 1.350 ;
        RECT  0.060 1.230 0.650 1.350 ;
    END
END AN3D0

MACRO AN3D1
    CLASS CORE ;
    FOREIGN AN3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.275 1.350 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.680 0.950 1.120 ;
        RECT  0.780 0.680 0.850 0.930 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.680 0.620 0.910 ;
        RECT  0.450 0.680 0.550 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.165 1.400 0.165 ;
        RECT  0.880 -0.165 1.070 0.300 ;
        RECT  0.000 -0.165 0.880 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.635 1.400 1.965 ;
        RECT  0.880 1.450 1.070 1.965 ;
        RECT  0.585 1.635 0.880 1.965 ;
        RECT  0.395 1.450 0.585 1.965 ;
        RECT  0.000 1.635 0.395 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.045 0.410 1.135 1.340 ;
        RECT  0.100 0.410 1.045 0.520 ;
        RECT  0.760 1.230 1.045 1.340 ;
        RECT  0.650 1.075 0.760 1.340 ;
        RECT  0.060 1.230 0.650 1.340 ;
    END
END AN3D1

MACRO AN3D2
    CLASS CORE ;
    FOREIGN AN3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.545 1.350 1.205 ;
        RECT  1.250 0.275 1.260 1.490 ;
        RECT  1.150 0.275 1.250 0.675 ;
        RECT  1.150 1.055 1.250 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.825 0.930 ;
        RECT  0.650 0.680 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.680 0.200 0.930 ;
        RECT  0.050 0.680 0.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 -0.165 1.600 0.165 ;
        RECT  1.405 -0.165 1.525 0.455 ;
        RECT  0.995 -0.165 1.405 0.165 ;
        RECT  0.845 -0.165 0.995 0.345 ;
        RECT  0.000 -0.165 0.845 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 1.635 1.600 1.965 ;
        RECT  1.405 1.325 1.525 1.965 ;
        RECT  0.770 1.635 1.405 1.965 ;
        RECT  0.770 1.390 1.040 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.315 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.035 0.775 1.140 0.945 ;
        RECT  0.935 0.450 1.035 1.300 ;
        RECT  0.060 0.450 0.935 0.560 ;
        RECT  0.205 1.210 0.935 1.300 ;
        RECT  0.085 1.210 0.205 1.450 ;
    END
END AN3D2

MACRO AN3D4
    CLASS CORE ;
    FOREIGN AN3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.310 2.505 0.690 ;
        RECT  2.450 1.110 2.505 1.490 ;
        RECT  2.150 0.310 2.450 1.490 ;
        RECT  1.850 0.310 2.150 0.690 ;
        RECT  1.850 1.110 2.150 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.730 1.580 0.940 ;
        RECT  1.450 0.500 1.550 0.940 ;
        RECT  0.360 0.500 1.450 0.590 ;
        RECT  0.270 0.500 0.360 0.780 ;
        RECT  0.190 0.680 0.270 0.780 ;
        RECT  0.050 0.680 0.190 1.120 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.220 0.700 1.350 1.100 ;
        RECT  0.550 1.010 1.220 1.100 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.700 0.950 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.735 -0.165 2.800 0.165 ;
        RECT  2.615 -0.165 2.735 0.690 ;
        RECT  0.180 -0.165 2.615 0.165 ;
        RECT  0.060 -0.165 0.180 0.570 ;
        RECT  0.000 -0.165 0.060 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.735 1.635 2.800 1.965 ;
        RECT  2.615 1.110 2.735 1.965 ;
        RECT  1.245 1.635 2.615 1.965 ;
        RECT  1.055 1.390 1.245 1.965 ;
        RECT  0.190 1.635 1.055 1.965 ;
        RECT  0.070 1.230 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.850 0.310 2.050 0.690 ;
        RECT  1.850 1.110 2.050 1.490 ;
        RECT  1.760 0.800 1.960 0.910 ;
        RECT  1.670 0.310 1.760 1.300 ;
        RECT  0.795 0.310 1.670 0.410 ;
        RECT  0.300 1.210 1.670 1.300 ;
    END
END AN3D4

MACRO AN3D8
    CLASS CORE ;
    FOREIGN AN3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.310 4.305 0.690 ;
        RECT  3.650 1.110 4.305 1.490 ;
        RECT  3.350 0.310 3.650 1.490 ;
        RECT  2.615 0.310 3.350 0.690 ;
        RECT  2.615 1.110 3.350 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.1645 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 0.710 2.300 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.555 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.750 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 -0.165 4.600 0.165 ;
        RECT  4.415 -0.165 4.535 0.690 ;
        RECT  2.045 -0.165 4.415 0.165 ;
        RECT  1.855 -0.165 2.045 0.410 ;
        RECT  0.000 -0.165 1.855 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 1.635 4.600 1.965 ;
        RECT  4.415 1.110 4.535 1.965 ;
        RECT  1.770 1.635 4.415 1.965 ;
        RECT  1.770 1.390 2.055 1.490 ;
        RECT  1.630 1.390 1.770 1.965 ;
        RECT  1.325 1.390 1.630 1.490 ;
        RECT  0.770 1.635 1.630 1.965 ;
        RECT  0.770 1.390 1.005 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.295 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 0.310 4.305 0.690 ;
        RECT  3.750 1.110 4.305 1.490 ;
        RECT  2.615 0.310 3.250 0.690 ;
        RECT  2.615 1.110 3.250 1.490 ;
        RECT  2.500 0.800 2.990 0.900 ;
        RECT  2.410 0.800 2.500 1.300 ;
        RECT  0.955 1.210 2.410 1.300 ;
        RECT  1.065 0.500 2.315 0.590 ;
        RECT  0.290 0.310 1.535 0.410 ;
        RECT  0.845 0.500 0.955 1.300 ;
        RECT  0.180 0.500 0.845 0.590 ;
        RECT  0.180 1.210 0.845 1.300 ;
        RECT  0.060 0.350 0.180 0.590 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AN3D8

MACRO AN3XD1
    CLASS CORE ;
    FOREIGN AN3XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.275 1.350 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.680 0.950 1.105 ;
        RECT  0.700 0.750 0.850 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.680 0.565 1.105 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.105 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.055 -0.165 1.400 0.165 ;
        RECT  0.865 -0.165 1.055 0.300 ;
        RECT  0.000 -0.165 0.865 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.635 1.400 1.965 ;
        RECT  0.770 1.395 1.090 1.485 ;
        RECT  0.630 1.395 0.770 1.965 ;
        RECT  0.285 1.395 0.630 1.485 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.045 0.410 1.135 1.305 ;
        RECT  0.045 0.410 1.045 0.520 ;
        RECT  0.175 1.215 1.045 1.305 ;
        RECT  0.085 1.215 0.175 1.460 ;
    END
END AN3XD1

MACRO AN4D0
    CLASS CORE ;
    FOREIGN AN4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.275 1.550 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.675 1.150 1.120 ;
        RECT  0.980 0.675 1.050 0.925 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.820 0.925 ;
        RECT  0.650 0.680 0.750 1.120 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.120 ;
        RECT  0.190 0.680 0.250 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.165 1.600 0.165 ;
        RECT  1.080 -0.165 1.270 0.300 ;
        RECT  0.000 -0.165 1.080 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.635 1.600 1.965 ;
        RECT  0.070 1.195 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.245 0.410 1.335 1.330 ;
        RECT  0.060 0.410 1.245 0.520 ;
        RECT  0.310 1.230 1.245 1.330 ;
    END
END AN4D0

MACRO AN4D1
    CLASS CORE ;
    FOREIGN AN4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.275 1.550 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0285 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.675 1.150 1.120 ;
        RECT  0.980 0.675 1.050 0.925 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.820 0.925 ;
        RECT  0.650 0.680 0.750 1.120 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.120 ;
        RECT  0.190 0.680 0.250 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.165 1.600 0.165 ;
        RECT  1.080 -0.165 1.270 0.300 ;
        RECT  0.000 -0.165 1.080 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.635 1.600 1.965 ;
        RECT  0.070 1.195 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.245 0.410 1.335 1.330 ;
        RECT  0.060 0.410 1.245 0.520 ;
        RECT  0.310 1.230 1.245 1.330 ;
    END
END AN4D1

MACRO AN4D2
    CLASS CORE ;
    FOREIGN AN4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.535 0.510 1.550 1.200 ;
        RECT  1.445 0.275 1.535 1.500 ;
        RECT  1.305 0.275 1.445 0.410 ;
        RECT  1.305 1.390 1.445 1.500 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  0.980 0.710 1.050 0.930 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.785 0.930 ;
        RECT  0.650 0.710 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.165 1.800 0.165 ;
        RECT  1.625 -0.165 1.735 0.445 ;
        RECT  0.000 -0.165 1.625 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 1.635 1.800 1.965 ;
        RECT  1.625 1.335 1.735 1.965 ;
        RECT  0.185 1.635 1.625 1.965 ;
        RECT  0.065 1.210 0.185 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.500 1.335 1.300 ;
        RECT  0.190 0.500 1.240 0.600 ;
        RECT  0.295 1.210 1.240 1.300 ;
        RECT  0.070 0.360 0.190 0.600 ;
    END
END AN4D2

MACRO AN4D4
    CLASS CORE ;
    FOREIGN AN4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.105 0.690 ;
        RECT  3.050 1.110 3.105 1.490 ;
        RECT  2.750 0.310 3.050 1.490 ;
        RECT  2.450 0.310 2.750 0.690 ;
        RECT  2.450 1.110 2.750 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.510 2.160 1.100 ;
        RECT  0.350 0.510 2.050 0.600 ;
        RECT  0.200 0.510 0.350 1.100 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 0.710 1.950 1.300 ;
        RECT  0.560 1.210 1.820 1.300 ;
        RECT  0.450 0.710 0.560 1.300 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.560 1.100 ;
        RECT  0.950 1.010 1.450 1.100 ;
        RECT  0.850 0.710 0.950 1.100 ;
        RECT  0.760 0.710 0.850 0.930 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.335 -0.165 3.400 0.165 ;
        RECT  3.215 -0.165 3.335 0.690 ;
        RECT  0.255 -0.165 3.215 0.165 ;
        RECT  0.075 -0.165 0.255 0.420 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.335 1.635 3.400 1.965 ;
        RECT  3.215 1.110 3.335 1.965 ;
        RECT  0.185 1.635 3.215 1.965 ;
        RECT  0.065 1.345 0.185 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.450 0.310 2.650 0.690 ;
        RECT  2.450 1.110 2.650 1.490 ;
        RECT  2.340 0.800 2.560 0.900 ;
        RECT  2.250 0.310 2.340 1.490 ;
        RECT  1.065 0.310 2.250 0.410 ;
        RECT  0.295 1.390 2.250 1.490 ;
    END
END AN4D4

MACRO AN4D8
    CLASS CORE ;
    FOREIGN AN4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.310 5.105 0.690 ;
        RECT  4.450 1.110 5.105 1.490 ;
        RECT  4.150 0.310 4.450 1.490 ;
        RECT  3.450 0.310 4.150 0.690 ;
        RECT  3.450 1.110 4.150 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.1645 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.710 3.005 0.890 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.710 2.405 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.195 0.710 1.605 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.195 0.710 0.605 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.335 -0.165 5.400 0.165 ;
        RECT  5.215 -0.165 5.335 0.690 ;
        RECT  2.970 -0.165 5.215 0.165 ;
        RECT  2.970 0.305 3.355 0.410 ;
        RECT  2.830 -0.165 2.970 0.410 ;
        RECT  0.000 -0.165 2.830 0.165 ;
        RECT  2.625 0.305 2.830 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.335 1.635 5.400 1.965 ;
        RECT  5.215 1.110 5.335 1.965 ;
        RECT  2.770 1.635 5.215 1.965 ;
        RECT  2.770 1.390 3.340 1.490 ;
        RECT  2.630 1.390 2.770 1.965 ;
        RECT  2.105 1.390 2.630 1.490 ;
        RECT  1.570 1.635 2.630 1.965 ;
        RECT  1.570 1.390 1.795 1.490 ;
        RECT  1.430 1.390 1.570 1.965 ;
        RECT  1.065 1.390 1.430 1.490 ;
        RECT  0.770 1.635 1.430 1.965 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.190 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        RECT  0.070 1.210 0.190 1.490 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.550 0.310 5.105 0.690 ;
        RECT  4.550 1.110 5.105 1.490 ;
        RECT  3.450 0.310 4.050 0.690 ;
        RECT  3.450 1.110 4.050 1.490 ;
        RECT  3.340 0.800 3.800 0.900 ;
        RECT  3.250 0.800 3.340 1.300 ;
        RECT  0.880 1.210 3.250 1.300 ;
        RECT  2.515 0.500 3.110 0.590 ;
        RECT  2.425 0.310 2.515 0.590 ;
        RECT  1.850 0.310 2.425 0.410 ;
        RECT  1.070 0.500 2.310 0.590 ;
        RECT  0.300 0.310 1.530 0.410 ;
        RECT  0.780 0.500 0.880 1.300 ;
        RECT  0.190 0.500 0.780 0.590 ;
        RECT  0.300 1.210 0.780 1.300 ;
        RECT  0.070 0.350 0.190 0.590 ;
    END
END AN4D8

MACRO AN4XD1
    CLASS CORE ;
    FOREIGN AN4XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.275 1.550 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.980 0.675 1.050 0.925 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.820 0.925 ;
        RECT  0.650 0.680 0.750 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.680 0.555 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.350 1.090 ;
        RECT  0.190 0.680 0.250 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.165 1.600 0.165 ;
        RECT  1.080 -0.165 1.270 0.300 ;
        RECT  0.000 -0.165 1.080 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.635 1.600 1.965 ;
        RECT  0.970 1.390 1.300 1.485 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.565 1.390 0.830 1.490 ;
        RECT  0.190 1.635 0.830 1.965 ;
        RECT  0.070 1.165 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.245 0.410 1.335 1.300 ;
        RECT  0.060 0.410 1.245 0.520 ;
        RECT  0.310 1.200 1.245 1.300 ;
    END
END AN4XD1

MACRO ANTENNA
    CLASS CORE ;
    FOREIGN ANTENNA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN I
        ANTENNADIFFAREA 0.1070 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.275 0.255 0.685 ;
        RECT  0.145 0.275 0.150 0.910 ;
        RECT  0.050 0.490 0.145 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 0.400 1.965 ;
        END
    END VDD
END ANTENNA

MACRO AO211D0
    CLASS CORE ;
    FOREIGN AO211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.285 1.550 1.490 ;
        RECT  1.365 0.285 1.450 0.410 ;
        RECT  1.405 1.065 1.450 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.970 0.700 1.050 0.950 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 -0.165 1.600 0.165 ;
        RECT  1.110 -0.165 1.240 0.410 ;
        RECT  0.670 -0.165 1.110 0.165 ;
        RECT  0.540 -0.165 0.670 0.410 ;
        RECT  0.000 -0.165 0.540 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.635 1.600 1.965 ;
        RECT  1.070 1.220 1.240 1.965 ;
        RECT  0.000 1.635 1.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.500 1.340 0.950 ;
        RECT  0.955 0.500 1.240 0.590 ;
        RECT  0.825 0.285 0.955 0.590 ;
        RECT  0.360 0.500 0.825 0.590 ;
        RECT  0.595 1.240 0.730 1.525 ;
        RECT  0.180 1.425 0.595 1.525 ;
        RECT  0.360 1.210 0.505 1.315 ;
        RECT  0.270 0.500 0.360 1.315 ;
        RECT  0.200 0.500 0.270 0.590 ;
        RECT  0.070 0.285 0.200 0.590 ;
        RECT  0.060 1.240 0.180 1.525 ;
    END
END AO211D0

MACRO AO211D1
    CLASS CORE ;
    FOREIGN AO211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.285 1.550 1.490 ;
        RECT  1.365 0.285 1.450 0.410 ;
        RECT  1.405 1.045 1.450 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.970 0.700 1.050 0.950 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 -0.165 1.600 0.165 ;
        RECT  1.100 -0.165 1.250 0.410 ;
        RECT  0.680 -0.165 1.100 0.165 ;
        RECT  0.530 -0.165 0.680 0.410 ;
        RECT  0.000 -0.165 0.530 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.635 1.600 1.965 ;
        RECT  1.110 1.210 1.240 1.965 ;
        RECT  0.000 1.635 1.110 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.500 1.340 0.940 ;
        RECT  0.360 0.500 1.240 0.590 ;
        RECT  0.610 1.240 0.730 1.510 ;
        RECT  0.180 1.410 0.610 1.510 ;
        RECT  0.360 1.210 0.495 1.300 ;
        RECT  0.270 0.500 0.360 1.300 ;
        RECT  0.180 0.500 0.270 0.590 ;
        RECT  0.060 0.350 0.180 0.590 ;
        RECT  0.060 1.240 0.180 1.510 ;
    END
END AO211D1

MACRO AO211D2
    CLASS CORE ;
    FOREIGN AO211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.505 1.550 1.300 ;
        RECT  1.300 0.505 1.450 0.655 ;
        RECT  1.300 1.200 1.450 1.300 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.500 1.150 0.900 ;
        RECT  0.955 0.725 1.050 0.900 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.815 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 -0.165 1.800 0.165 ;
        RECT  1.170 0.310 1.740 0.410 ;
        RECT  1.030 -0.165 1.170 0.410 ;
        RECT  0.000 -0.165 1.030 0.165 ;
        RECT  0.480 0.310 1.030 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.635 1.800 1.965 ;
        RECT  1.370 1.390 1.740 1.490 ;
        RECT  1.230 1.390 1.370 1.965 ;
        RECT  1.010 1.390 1.230 1.490 ;
        RECT  0.000 1.635 1.230 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.765 1.340 1.110 ;
        RECT  1.155 1.010 1.240 1.110 ;
        RECT  1.055 1.010 1.155 1.300 ;
        RECT  0.360 1.210 1.055 1.300 ;
        RECT  0.360 0.500 0.940 0.590 ;
        RECT  0.060 1.390 0.770 1.515 ;
        RECT  0.270 0.500 0.360 1.300 ;
        RECT  0.185 0.500 0.270 0.590 ;
        RECT  0.065 0.350 0.185 0.590 ;
    END
END AO211D2

MACRO AO211D4
    CLASS CORE ;
    FOREIGN AO211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.310 3.305 0.690 ;
        RECT  3.250 1.110 3.305 1.490 ;
        RECT  2.950 0.310 3.250 1.490 ;
        RECT  2.650 0.310 2.950 0.690 ;
        RECT  2.650 1.110 2.950 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.700 1.150 1.100 ;
        RECT  0.190 1.010 1.010 1.100 ;
        RECT  0.050 0.700 0.190 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.700 2.150 1.100 ;
        RECT  1.390 1.010 2.050 1.100 ;
        RECT  1.250 0.700 1.390 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.950 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 -0.165 3.600 0.165 ;
        RECT  3.415 -0.165 3.535 0.705 ;
        RECT  1.170 -0.165 3.415 0.165 ;
        RECT  1.170 0.310 2.320 0.410 ;
        RECT  1.030 -0.165 1.170 0.410 ;
        RECT  0.000 -0.165 1.030 0.165 ;
        RECT  0.190 0.310 1.030 0.410 ;
        RECT  0.070 0.310 0.190 0.570 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 1.635 3.600 1.965 ;
        RECT  3.415 1.095 3.535 1.965 ;
        RECT  0.750 1.635 3.415 1.965 ;
        RECT  0.560 1.390 0.750 1.965 ;
        RECT  0.000 1.635 0.560 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.650 0.310 2.850 0.690 ;
        RECT  2.650 1.110 2.850 1.490 ;
        RECT  2.395 0.800 2.760 0.900 ;
        RECT  2.305 0.500 2.395 1.300 ;
        RECT  1.225 1.390 2.320 1.490 ;
        RECT  0.300 0.500 2.305 0.590 ;
        RECT  1.340 1.210 2.305 1.300 ;
        RECT  1.110 1.210 1.225 1.490 ;
        RECT  0.200 1.210 1.110 1.300 ;
        RECT  0.065 1.210 0.200 1.450 ;
    END
END AO211D4

MACRO AO21D0
    CLASS CORE ;
    FOREIGN AO21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.275 1.350 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.680 0.790 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.165 1.400 0.165 ;
        RECT  0.880 -0.165 1.030 0.370 ;
        RECT  0.180 -0.165 0.880 0.165 ;
        RECT  0.070 -0.165 0.180 0.475 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.635 1.400 1.965 ;
        RECT  0.880 1.240 1.030 1.965 ;
        RECT  0.000 1.635 0.880 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.460 1.105 0.940 ;
        RECT  0.725 0.460 0.990 0.560 ;
        RECT  0.595 0.275 0.725 0.560 ;
        RECT  0.595 1.240 0.725 1.525 ;
        RECT  0.360 0.470 0.595 0.560 ;
        RECT  0.180 1.425 0.595 1.525 ;
        RECT  0.360 1.210 0.485 1.300 ;
        RECT  0.270 0.470 0.360 1.300 ;
        RECT  0.070 1.240 0.180 1.525 ;
    END
END AO21D0

MACRO AO21D1
    CLASS CORE ;
    FOREIGN AO21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.275 1.350 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.810 0.950 ;
        RECT  0.650 0.680 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.165 1.400 0.165 ;
        RECT  0.880 -0.165 1.030 0.370 ;
        RECT  0.190 -0.165 0.880 0.165 ;
        RECT  0.070 -0.165 0.190 0.570 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.635 1.400 1.965 ;
        RECT  0.880 1.410 1.030 1.965 ;
        RECT  0.000 1.635 0.880 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.005 0.460 1.105 1.300 ;
        RECT  0.555 0.460 1.005 0.560 ;
        RECT  0.305 1.210 1.005 1.300 ;
        RECT  0.190 1.390 0.765 1.490 ;
        RECT  0.070 1.240 0.190 1.490 ;
    END
END AO21D1

MACRO AO21D2
    CLASS CORE ;
    FOREIGN AO21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.545 1.350 1.195 ;
        RECT  1.250 0.275 1.260 1.490 ;
        RECT  1.160 0.275 1.250 0.675 ;
        RECT  1.160 1.045 1.250 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.810 0.950 ;
        RECT  0.650 0.680 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.530 -0.165 1.600 0.165 ;
        RECT  1.410 -0.165 1.530 0.465 ;
        RECT  1.000 -0.165 1.410 0.165 ;
        RECT  0.850 -0.165 1.000 0.370 ;
        RECT  0.190 -0.165 0.850 0.165 ;
        RECT  0.070 -0.165 0.190 0.570 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.530 1.635 1.600 1.965 ;
        RECT  1.410 1.325 1.530 1.965 ;
        RECT  1.045 1.635 1.410 1.965 ;
        RECT  0.855 1.390 1.045 1.965 ;
        RECT  0.000 1.635 0.855 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.460 1.050 1.300 ;
        RECT  0.535 0.460 0.950 0.560 ;
        RECT  0.305 1.210 0.950 1.300 ;
        RECT  0.190 1.390 0.745 1.490 ;
        RECT  0.070 1.240 0.190 1.490 ;
    END
END AO21D2

MACRO AO21D4
    CLASS CORE ;
    FOREIGN AO21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.310 2.550 0.690 ;
        RECT  2.450 1.110 2.550 1.490 ;
        RECT  2.150 0.310 2.450 1.490 ;
        RECT  1.870 0.310 2.150 0.690 ;
        RECT  1.870 1.110 2.150 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.730 1.580 0.940 ;
        RECT  1.450 0.500 1.550 0.940 ;
        RECT  0.170 0.500 1.450 0.590 ;
        RECT  0.050 0.500 0.170 1.120 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.700 0.950 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.700 1.350 1.100 ;
        RECT  0.550 1.010 1.240 1.100 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.870 0.310 2.050 0.690 ;
        RECT  1.870 1.110 2.050 1.490 ;
        RECT  1.760 0.800 1.970 0.900 ;
        RECT  1.670 0.310 1.760 1.300 ;
        RECT  0.275 0.310 1.670 0.410 ;
        RECT  0.535 1.210 1.670 1.300 ;
        RECT  0.275 1.390 1.525 1.490 ;
    END
END AO21D4

MACRO AO221D0
    CLASS CORE ;
    FOREIGN AO221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.825 0.285 1.950 1.290 ;
        RECT  1.810 0.285 1.825 0.455 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.710 1.550 1.105 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.895 0.530 1.065 0.640 ;
        RECT  0.160 0.530 0.895 0.620 ;
        RECT  0.050 0.530 0.160 1.235 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.350 1.090 ;
        RECT  1.075 0.800 1.245 0.930 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.780 0.970 1.090 ;
        RECT  0.775 0.780 0.845 0.915 ;
        RECT  0.640 0.710 0.775 0.915 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.375 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.695 1.635 2.000 1.965 ;
        RECT  1.525 1.445 1.695 1.965 ;
        RECT  0.000 1.635 1.525 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.720 0.530 1.735 1.305 ;
        RECT  1.640 0.310 1.720 1.305 ;
        RECT  1.620 0.310 1.640 0.620 ;
        RECT  0.710 1.215 1.640 1.305 ;
        RECT  0.255 0.310 1.620 0.420 ;
        RECT  0.210 1.415 1.365 1.525 ;
        RECT  0.580 1.030 0.710 1.305 ;
        RECT  0.080 1.345 0.210 1.525 ;
    END
END AO221D0

MACRO AO221D1
    CLASS CORE ;
    FOREIGN AO221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.285 2.150 1.490 ;
        RECT  1.965 0.285 2.050 0.410 ;
        RECT  2.005 1.045 2.050 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.750 1.100 ;
        RECT  1.580 0.700 1.650 0.950 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.700 1.150 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.700 1.410 0.950 ;
        RECT  1.250 0.700 1.350 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.190 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.700 0.755 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.850 -0.165 2.200 0.165 ;
        RECT  1.700 -0.165 1.850 0.410 ;
        RECT  1.040 -0.165 1.700 0.165 ;
        RECT  0.890 -0.165 1.040 0.410 ;
        RECT  0.225 -0.165 0.890 0.165 ;
        RECT  0.105 -0.165 0.225 0.565 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.635 2.200 1.965 ;
        RECT  1.705 1.210 1.840 1.965 ;
        RECT  0.000 1.635 1.705 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 0.500 1.940 0.950 ;
        RECT  0.435 0.500 1.840 0.590 ;
        RECT  0.870 1.390 1.595 1.490 ;
        RECT  0.755 1.210 1.335 1.300 ;
        RECT  0.640 1.210 0.755 1.500 ;
        RECT  0.075 1.390 0.640 1.500 ;
        RECT  0.435 1.160 0.530 1.280 ;
        RECT  0.335 0.500 0.435 1.280 ;
    END
END AO221D1

MACRO AO221D2
    CLASS CORE ;
    FOREIGN AO221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.535 2.150 1.195 ;
        RECT  2.050 0.275 2.065 1.490 ;
        RECT  1.955 0.275 2.050 0.675 ;
        RECT  1.955 1.045 2.050 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.630 0.950 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.700 1.010 0.950 ;
        RECT  0.850 0.700 0.950 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.165 2.400 0.165 ;
        RECT  2.210 -0.165 2.330 0.455 ;
        RECT  1.370 -0.165 2.210 0.165 ;
        RECT  1.370 0.320 1.830 0.410 ;
        RECT  1.230 -0.165 1.370 0.410 ;
        RECT  0.225 -0.165 1.230 0.165 ;
        RECT  0.840 0.320 1.230 0.410 ;
        RECT  0.105 -0.165 0.225 0.590 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.635 2.400 1.965 ;
        RECT  2.210 1.325 2.330 1.965 ;
        RECT  1.810 1.635 2.210 1.965 ;
        RECT  1.695 1.095 1.810 1.965 ;
        RECT  0.000 1.635 1.695 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 0.775 1.910 0.945 ;
        RECT  1.740 0.500 1.840 0.945 ;
        RECT  0.435 0.500 1.740 0.590 ;
        RECT  0.875 1.390 1.585 1.490 ;
        RECT  0.740 1.210 1.325 1.300 ;
        RECT  0.640 1.210 0.740 1.500 ;
        RECT  0.075 1.390 0.640 1.500 ;
        RECT  0.435 1.170 0.525 1.280 ;
        RECT  0.335 0.500 0.435 1.280 ;
    END
END AO221D2

MACRO AO221D4
    CLASS CORE ;
    FOREIGN AO221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.310 4.105 0.690 ;
        RECT  4.050 1.110 4.105 1.490 ;
        RECT  3.750 0.310 4.050 1.490 ;
        RECT  3.450 0.310 3.750 0.690 ;
        RECT  3.450 1.110 3.750 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.700 0.360 1.100 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.350 0.900 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.750 1.100 ;
        RECT  0.950 1.010 1.650 1.100 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.765 0.700 0.850 0.920 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.700 2.750 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.700 2.950 1.100 ;
        RECT  2.150 1.010 2.850 1.100 ;
        RECT  2.040 0.700 2.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.335 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.335 0.690 ;
        RECT  2.610 -0.165 4.215 0.165 ;
        RECT  2.420 -0.165 2.610 0.410 ;
        RECT  0.770 -0.165 2.420 0.165 ;
        RECT  0.770 0.310 1.280 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.295 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.335 1.635 4.400 1.965 ;
        RECT  4.215 1.110 4.335 1.965 ;
        RECT  0.490 1.635 4.215 1.965 ;
        RECT  0.300 1.390 0.490 1.965 ;
        RECT  0.000 1.635 0.300 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.450 0.310 3.650 0.690 ;
        RECT  3.450 1.110 3.650 1.490 ;
        RECT  3.215 0.800 3.560 0.900 ;
        RECT  3.105 0.500 3.215 1.300 ;
        RECT  0.185 0.500 3.105 0.590 ;
        RECT  1.900 1.210 3.105 1.300 ;
        RECT  0.810 1.390 2.880 1.490 ;
        RECT  0.185 1.210 1.790 1.300 ;
        RECT  0.065 0.350 0.185 0.590 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AO221D4

MACRO AO222D0
    CLASS CORE ;
    FOREIGN AO222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.225 0.300 2.350 1.290 ;
        RECT  2.145 0.300 2.225 0.415 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.710 1.950 1.090 ;
        RECT  1.650 0.755 1.840 0.925 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.510 1.555 0.915 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0285 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 0.530 1.035 0.640 ;
        RECT  0.160 0.530 0.865 0.620 ;
        RECT  0.050 0.530 0.160 1.235 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.350 1.090 ;
        RECT  1.040 0.800 1.245 0.930 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.780 0.950 1.090 ;
        RECT  0.775 0.780 0.845 0.915 ;
        RECT  0.640 0.710 0.775 0.915 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.375 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 -0.165 2.400 0.165 ;
        RECT  1.845 -0.165 2.030 0.420 ;
        RECT  0.000 -0.165 1.845 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.150 1.635 2.400 1.965 ;
        RECT  1.980 1.445 2.150 1.965 ;
        RECT  0.000 1.635 1.980 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.040 0.510 2.135 1.305 ;
        RECT  1.755 0.510 2.040 0.600 ;
        RECT  0.710 1.215 2.040 1.305 ;
        RECT  0.210 1.415 1.870 1.525 ;
        RECT  1.665 0.310 1.755 0.600 ;
        RECT  0.255 0.310 1.665 0.420 ;
        RECT  0.580 1.030 0.710 1.305 ;
        RECT  0.080 1.345 0.210 1.525 ;
    END
END AO222D0

MACRO AO222D1
    CLASS CORE ;
    FOREIGN AO222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.275 2.350 1.490 ;
        RECT  2.210 0.275 2.250 0.675 ;
        RECT  2.210 1.045 2.250 1.490 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.700 1.880 0.950 ;
        RECT  1.650 0.700 1.750 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.155 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.165 2.400 0.165 ;
        RECT  1.900 -0.165 2.050 0.390 ;
        RECT  0.770 -0.165 1.900 0.165 ;
        RECT  0.770 0.300 1.290 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.060 0.300 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.065 1.635 2.400 1.965 ;
        RECT  1.950 1.100 2.065 1.965 ;
        RECT  1.385 1.390 1.950 1.490 ;
        RECT  0.000 1.635 1.950 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.100 0.760 2.140 0.930 ;
        RECT  2.000 0.500 2.100 0.930 ;
        RECT  0.350 0.500 2.000 0.590 ;
        RECT  0.820 1.210 1.840 1.300 ;
        RECT  0.060 1.390 1.270 1.500 ;
        RECT  0.350 1.210 0.500 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
    END
END AO222D1

MACRO AO222D2
    CLASS CORE ;
    FOREIGN AO222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.260 0.535 2.350 1.195 ;
        RECT  2.250 0.275 2.260 1.490 ;
        RECT  2.160 0.275 2.250 0.675 ;
        RECT  2.160 1.045 2.250 1.490 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.700 1.830 0.950 ;
        RECT  1.650 0.700 1.750 1.090 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.090 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.155 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.800 0.950 ;
        RECT  0.650 0.700 0.750 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.165 2.600 0.165 ;
        RECT  2.410 -0.165 2.530 0.455 ;
        RECT  2.000 -0.165 2.410 0.165 ;
        RECT  1.850 -0.165 2.000 0.390 ;
        RECT  0.770 -0.165 1.850 0.165 ;
        RECT  0.770 0.300 1.255 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.060 0.300 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 1.635 2.600 1.965 ;
        RECT  2.410 1.325 2.530 1.965 ;
        RECT  1.770 1.635 2.410 1.965 ;
        RECT  1.770 1.380 2.045 1.500 ;
        RECT  1.630 1.380 1.770 1.965 ;
        RECT  1.345 1.380 1.630 1.500 ;
        RECT  0.000 1.635 1.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.050 0.760 2.090 0.930 ;
        RECT  1.950 0.500 2.050 0.930 ;
        RECT  0.360 0.500 1.950 0.590 ;
        RECT  0.815 1.200 1.795 1.290 ;
        RECT  0.700 1.380 1.255 1.500 ;
        RECT  0.600 1.230 0.700 1.500 ;
        RECT  0.180 1.400 0.600 1.500 ;
        RECT  0.360 1.200 0.485 1.290 ;
        RECT  0.270 0.500 0.360 1.290 ;
        RECT  0.060 1.230 0.180 1.500 ;
    END
END AO222D2

MACRO AO222D4
    CLASS CORE ;
    FOREIGN AO222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.430 4.685 0.620 ;
        RECT  4.450 1.105 4.685 1.295 ;
        RECT  4.150 0.430 4.450 1.295 ;
        RECT  3.965 0.430 4.150 0.620 ;
        RECT  3.965 1.105 4.150 1.295 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.700 1.150 1.100 ;
        RECT  0.170 1.010 1.030 1.100 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.700 2.150 1.100 ;
        RECT  1.370 1.010 2.050 1.100 ;
        RECT  1.250 0.700 1.370 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.950 0.900 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.700 3.150 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.700 3.400 0.920 ;
        RECT  3.250 0.700 3.350 1.100 ;
        RECT  2.750 1.010 3.250 1.100 ;
        RECT  2.650 0.700 2.750 1.100 ;
        RECT  2.450 0.700 2.650 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 -0.165 5.000 0.165 ;
        RECT  4.810 -0.165 4.930 0.685 ;
        RECT  4.420 -0.165 4.810 0.165 ;
        RECT  4.230 -0.165 4.420 0.325 ;
        RECT  3.830 -0.165 4.230 0.165 ;
        RECT  3.730 -0.165 3.830 0.685 ;
        RECT  2.570 -0.165 3.730 0.165 ;
        RECT  2.570 0.310 3.105 0.410 ;
        RECT  2.430 -0.165 2.570 0.410 ;
        RECT  0.770 -0.165 2.430 0.165 ;
        RECT  2.105 0.310 2.430 0.410 ;
        RECT  0.770 0.310 1.275 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.190 0.310 0.630 0.410 ;
        RECT  0.070 0.310 0.190 0.570 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 1.635 5.000 1.965 ;
        RECT  4.810 1.105 4.930 1.965 ;
        RECT  4.410 1.635 4.810 1.965 ;
        RECT  4.240 1.415 4.410 1.965 ;
        RECT  3.830 1.635 4.240 1.965 ;
        RECT  3.730 1.105 3.830 1.965 ;
        RECT  0.770 1.635 3.730 1.965 ;
        RECT  0.770 1.390 1.015 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.290 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.550 0.430 4.685 0.620 ;
        RECT  4.550 1.105 4.685 1.295 ;
        RECT  3.965 0.430 4.050 0.620 ;
        RECT  3.965 1.105 4.050 1.295 ;
        RECT  3.620 0.780 4.040 0.890 ;
        RECT  3.530 0.500 3.620 1.300 ;
        RECT  0.555 0.500 3.530 0.590 ;
        RECT  2.550 1.210 3.530 1.300 ;
        RECT  1.325 1.390 3.365 1.490 ;
        RECT  2.430 1.060 2.550 1.300 ;
        RECT  0.180 1.210 2.315 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO222D4

MACRO AO22D0
    CLASS CORE ;
    FOREIGN AO22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0830 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.310 1.550 1.490 ;
        RECT  1.340 0.310 1.440 0.425 ;
        RECT  1.360 1.365 1.440 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.555 0.170 0.745 ;
        RECT  0.050 0.555 0.150 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.710 1.170 1.090 ;
        RECT  1.010 0.710 1.030 0.835 ;
        RECT  0.900 0.490 1.010 0.835 ;
        RECT  0.560 0.490 0.900 0.585 ;
        RECT  0.430 0.490 0.560 0.690 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 0.965 0.860 1.090 ;
        RECT  0.650 0.680 0.760 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.555 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.165 1.600 0.165 ;
        RECT  0.065 -0.165 0.195 0.445 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.635 1.600 1.965 ;
        RECT  1.100 1.365 1.270 1.965 ;
        RECT  0.195 1.635 1.100 1.965 ;
        RECT  0.075 1.235 0.195 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.515 1.350 1.275 ;
        RECT  1.230 0.515 1.260 0.605 ;
        RECT  0.750 1.185 1.260 1.275 ;
        RECT  1.120 0.290 1.230 0.605 ;
        RECT  0.485 0.290 1.120 0.400 ;
        RECT  0.840 1.365 1.010 1.525 ;
        RECT  0.455 1.435 0.840 1.525 ;
        RECT  0.580 1.185 0.750 1.345 ;
        RECT  0.325 1.260 0.455 1.525 ;
    END
END AO22D0

MACRO AO22D1
    CLASS CORE ;
    FOREIGN AO22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.275 1.750 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.810 0.950 ;
        RECT  0.650 0.680 0.750 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.680 1.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 -0.165 1.800 0.165 ;
        RECT  0.580 -0.165 0.750 0.345 ;
        RECT  0.000 -0.165 0.580 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 1.635 1.800 1.965 ;
        RECT  0.310 1.390 0.500 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.345 0.450 1.460 1.300 ;
        RECT  0.060 0.450 1.345 0.560 ;
        RECT  0.830 1.210 1.345 1.300 ;
        RECT  0.715 1.390 1.290 1.490 ;
        RECT  0.615 1.210 0.715 1.490 ;
        RECT  0.195 1.210 0.615 1.300 ;
        RECT  0.075 1.210 0.195 1.450 ;
    END
END AO22D1

MACRO AO22D2
    CLASS CORE ;
    FOREIGN AO22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.860 0.535 1.950 1.195 ;
        RECT  1.850 0.275 1.860 1.490 ;
        RECT  1.760 0.275 1.850 0.675 ;
        RECT  1.760 1.045 1.850 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.810 0.950 ;
        RECT  0.650 0.680 0.750 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.680 1.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 -0.165 2.200 0.165 ;
        RECT  2.010 -0.165 2.130 0.455 ;
        RECT  1.610 -0.165 2.010 0.165 ;
        RECT  1.440 -0.165 1.610 0.345 ;
        RECT  0.750 -0.165 1.440 0.165 ;
        RECT  0.580 -0.165 0.750 0.345 ;
        RECT  0.000 -0.165 0.580 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 1.635 2.200 1.965 ;
        RECT  2.010 1.325 2.130 1.965 ;
        RECT  1.610 1.635 2.010 1.965 ;
        RECT  1.440 1.420 1.610 1.965 ;
        RECT  0.500 1.635 1.440 1.965 ;
        RECT  0.310 1.390 0.500 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.500 0.450 1.600 1.300 ;
        RECT  0.060 0.450 1.500 0.560 ;
        RECT  0.830 1.210 1.500 1.300 ;
        RECT  0.715 1.390 1.290 1.490 ;
        RECT  0.615 1.210 0.715 1.490 ;
        RECT  0.195 1.210 0.615 1.300 ;
        RECT  0.075 1.210 0.195 1.450 ;
    END
END AO22D2

MACRO AO22D4
    CLASS CORE ;
    FOREIGN AO22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.310 3.305 0.690 ;
        RECT  3.250 1.110 3.305 1.490 ;
        RECT  2.950 0.310 3.250 1.490 ;
        RECT  2.650 0.310 2.950 0.690 ;
        RECT  2.650 1.110 2.950 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.700 1.150 1.100 ;
        RECT  0.180 1.010 1.020 1.100 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.700 2.150 1.100 ;
        RECT  1.370 1.010 2.050 1.100 ;
        RECT  1.250 0.700 1.370 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.950 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 -0.165 3.600 0.165 ;
        RECT  3.415 -0.165 3.535 0.690 ;
        RECT  1.170 -0.165 3.415 0.165 ;
        RECT  1.170 0.310 2.320 0.410 ;
        RECT  1.030 -0.165 1.170 0.410 ;
        RECT  0.000 -0.165 1.030 0.165 ;
        RECT  0.180 0.310 1.030 0.410 ;
        RECT  0.060 0.310 0.180 0.560 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 1.635 3.600 1.965 ;
        RECT  3.415 1.110 3.535 1.965 ;
        RECT  0.770 1.635 3.415 1.965 ;
        RECT  0.770 1.390 1.015 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.295 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.650 0.310 2.850 0.690 ;
        RECT  2.650 1.110 2.850 1.490 ;
        RECT  2.405 0.800 2.765 0.900 ;
        RECT  2.290 0.500 2.405 1.300 ;
        RECT  1.225 1.390 2.320 1.490 ;
        RECT  0.550 0.500 2.290 0.590 ;
        RECT  1.340 1.210 2.290 1.300 ;
        RECT  1.125 1.210 1.225 1.490 ;
        RECT  0.185 1.210 1.125 1.300 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AO22D4

MACRO AO31D0
    CLASS CORE ;
    FOREIGN AO31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.285 1.550 1.490 ;
        RECT  1.395 0.285 1.450 0.480 ;
        RECT  1.425 1.255 1.450 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.910 1.170 1.290 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.550 1.165 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.930 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 -0.165 1.600 0.165 ;
        RECT  1.090 -0.165 1.260 0.400 ;
        RECT  0.235 -0.165 1.090 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 1.635 1.600 1.965 ;
        RECT  1.125 1.390 1.305 1.965 ;
        RECT  0.000 1.635 1.125 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.620 1.350 0.800 ;
        RECT  1.170 0.510 1.260 0.800 ;
        RECT  0.955 0.510 1.170 0.600 ;
        RECT  0.825 0.285 0.955 0.600 ;
        RECT  0.350 0.510 0.825 0.600 ;
        RECT  0.640 1.075 0.760 1.375 ;
        RECT  0.350 1.275 0.640 1.375 ;
        RECT  0.260 0.510 0.350 1.375 ;
        RECT  0.190 1.275 0.260 1.375 ;
        RECT  0.065 1.275 0.190 1.490 ;
    END
END AO31D0

MACRO AO31D1
    CLASS CORE ;
    FOREIGN AO31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.285 1.550 1.490 ;
        RECT  1.365 0.285 1.450 0.410 ;
        RECT  1.405 1.045 1.450 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 -0.165 1.600 0.165 ;
        RECT  1.100 -0.165 1.250 0.390 ;
        RECT  0.235 -0.165 1.100 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 1.635 1.600 1.965 ;
        RECT  1.125 1.245 1.265 1.965 ;
        RECT  0.000 1.635 1.125 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.500 1.340 0.930 ;
        RECT  0.350 0.500 1.240 0.590 ;
        RECT  0.295 1.390 1.015 1.490 ;
        RECT  0.350 1.210 0.760 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 1.210 0.260 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO31D1

MACRO AO31D2
    CLASS CORE ;
    FOREIGN AO31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.535 0.575 1.550 1.185 ;
        RECT  1.475 0.300 1.535 1.185 ;
        RECT  1.450 0.300 1.475 1.490 ;
        RECT  1.445 0.300 1.450 0.675 ;
        RECT  1.345 1.045 1.450 1.490 ;
        RECT  1.325 0.300 1.445 0.410 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.165 1.800 0.165 ;
        RECT  1.625 -0.165 1.735 0.465 ;
        RECT  1.235 -0.165 1.625 0.165 ;
        RECT  1.055 -0.165 1.235 0.410 ;
        RECT  0.235 -0.165 1.055 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 1.635 1.800 1.965 ;
        RECT  1.605 1.295 1.735 1.965 ;
        RECT  0.000 1.635 1.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.500 1.335 0.930 ;
        RECT  0.350 0.500 1.240 0.590 ;
        RECT  0.290 1.390 1.015 1.490 ;
        RECT  0.350 1.210 0.755 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 1.210 0.260 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO31D2

MACRO AO31D4
    CLASS CORE ;
    FOREIGN AO31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.310 3.305 0.690 ;
        RECT  3.250 1.110 3.305 1.490 ;
        RECT  2.950 0.310 3.250 1.490 ;
        RECT  2.650 0.310 2.950 0.690 ;
        RECT  2.650 1.110 2.950 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.700 2.150 0.900 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.780 1.695 0.890 ;
        RECT  1.450 0.500 1.550 0.890 ;
        RECT  0.360 0.500 1.450 0.590 ;
        RECT  0.270 0.500 0.360 0.780 ;
        RECT  0.170 0.680 0.270 0.780 ;
        RECT  0.050 0.680 0.170 1.120 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.350 1.100 ;
        RECT  0.550 1.010 1.250 1.100 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.700 0.950 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 -0.165 3.600 0.165 ;
        RECT  3.415 -0.165 3.535 0.690 ;
        RECT  2.320 -0.165 3.415 0.165 ;
        RECT  2.130 -0.165 2.320 0.410 ;
        RECT  0.180 -0.165 2.130 0.165 ;
        RECT  0.060 -0.165 0.180 0.570 ;
        RECT  0.000 -0.165 0.060 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 1.635 3.600 1.965 ;
        RECT  3.415 1.110 3.535 1.965 ;
        RECT  2.060 1.635 3.415 1.965 ;
        RECT  1.870 1.390 2.060 1.965 ;
        RECT  0.000 1.635 1.870 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.650 0.310 2.850 0.690 ;
        RECT  2.650 1.110 2.850 1.490 ;
        RECT  2.405 0.800 2.760 0.900 ;
        RECT  2.305 0.500 2.405 1.100 ;
        RECT  1.755 1.210 2.320 1.300 ;
        RECT  2.015 0.500 2.305 0.590 ;
        RECT  1.550 1.010 2.305 1.100 ;
        RECT  1.915 0.310 2.015 0.590 ;
        RECT  0.810 0.310 1.915 0.410 ;
        RECT  1.655 1.210 1.755 1.490 ;
        RECT  0.195 1.390 1.655 1.490 ;
        RECT  1.450 1.010 1.550 1.300 ;
        RECT  0.310 1.210 1.450 1.300 ;
        RECT  0.075 1.240 0.195 1.490 ;
    END
END AO31D4

MACRO AO32D0
    CLASS CORE ;
    FOREIGN AO32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.275 2.150 1.490 ;
        RECT  1.975 0.275 2.050 0.480 ;
        RECT  1.975 1.225 2.050 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.395 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.090 ;
        RECT  1.000 0.700 1.050 0.950 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.700 0.830 0.950 ;
        RECT  0.645 0.700 0.755 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.165 2.200 0.165 ;
        RECT  1.370 0.310 1.865 0.410 ;
        RECT  1.230 -0.165 1.370 0.410 ;
        RECT  0.235 -0.165 1.230 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.830 1.635 2.200 1.965 ;
        RECT  1.690 1.225 1.830 1.965 ;
        RECT  0.000 1.635 1.690 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.745 0.500 1.875 0.950 ;
        RECT  1.010 0.500 1.745 0.590 ;
        RECT  1.415 1.210 1.545 1.460 ;
        RECT  1.015 1.210 1.415 1.300 ;
        RECT  0.905 1.210 1.015 1.525 ;
        RECT  0.870 0.275 1.010 0.590 ;
        RECT  0.310 1.435 0.905 1.525 ;
        RECT  0.350 0.500 0.870 0.590 ;
        RECT  0.350 1.210 0.795 1.345 ;
        RECT  0.260 0.500 0.350 1.345 ;
        RECT  0.185 1.210 0.260 1.345 ;
        RECT  0.075 1.210 0.185 1.490 ;
    END
END AO32D0

MACRO AO32D1
    CLASS CORE ;
    FOREIGN AO32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.015 0.275 2.150 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.165 2.200 0.165 ;
        RECT  1.770 0.310 1.905 0.410 ;
        RECT  1.630 -0.165 1.770 0.410 ;
        RECT  0.235 -0.165 1.630 0.165 ;
        RECT  1.290 0.310 1.630 0.410 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.635 2.200 1.965 ;
        RECT  1.735 1.085 1.870 1.965 ;
        RECT  1.265 1.635 1.735 1.965 ;
        RECT  1.075 1.390 1.265 1.965 ;
        RECT  0.000 1.635 1.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.800 0.500 1.900 0.950 ;
        RECT  0.350 0.500 1.800 0.590 ;
        RECT  0.960 1.210 1.525 1.300 ;
        RECT  0.860 1.210 0.960 1.490 ;
        RECT  0.295 1.390 0.860 1.490 ;
        RECT  0.350 1.210 0.745 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 1.210 0.260 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO32D1

MACRO AO32D2
    CLASS CORE ;
    FOREIGN AO32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.535 2.150 1.195 ;
        RECT  2.050 0.275 2.060 1.490 ;
        RECT  1.960 0.275 2.050 0.675 ;
        RECT  1.960 1.045 2.050 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.165 2.400 0.165 ;
        RECT  2.210 -0.165 2.330 0.455 ;
        RECT  1.570 -0.165 2.210 0.165 ;
        RECT  1.570 0.310 1.850 0.410 ;
        RECT  1.430 -0.165 1.570 0.410 ;
        RECT  0.235 -0.165 1.430 0.165 ;
        RECT  1.285 0.310 1.430 0.410 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.635 2.400 1.965 ;
        RECT  2.210 1.345 2.330 1.965 ;
        RECT  1.815 1.635 2.210 1.965 ;
        RECT  1.685 1.080 1.815 1.965 ;
        RECT  1.265 1.635 1.685 1.965 ;
        RECT  1.075 1.390 1.265 1.965 ;
        RECT  0.000 1.635 1.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.750 0.500 1.850 0.930 ;
        RECT  0.350 0.500 1.750 0.590 ;
        RECT  0.960 1.210 1.525 1.300 ;
        RECT  0.860 1.210 0.960 1.490 ;
        RECT  0.295 1.390 0.860 1.490 ;
        RECT  0.350 1.210 0.745 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 1.210 0.260 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO32D2

MACRO AO32D4
    CLASS CORE ;
    FOREIGN AO32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.510 3.895 0.675 ;
        RECT  3.650 1.110 3.895 1.290 ;
        RECT  3.350 0.510 3.650 1.290 ;
        RECT  3.195 0.510 3.350 0.675 ;
        RECT  3.195 1.110 3.350 1.290 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.700 1.065 0.920 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.170 1.010 0.850 1.100 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.700 2.645 0.900 ;
        RECT  2.450 0.500 2.550 0.900 ;
        RECT  1.750 0.500 2.450 0.590 ;
        RECT  1.650 0.500 1.750 0.660 ;
        RECT  1.350 0.570 1.650 0.660 ;
        RECT  1.235 0.570 1.350 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.700 2.360 1.100 ;
        RECT  1.575 1.010 2.250 1.100 ;
        RECT  1.450 0.775 1.575 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.700 2.150 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.005 -0.165 4.125 0.675 ;
        RECT  3.640 -0.165 4.005 0.165 ;
        RECT  3.450 -0.165 3.640 0.410 ;
        RECT  3.050 -0.165 3.450 0.165 ;
        RECT  2.860 -0.165 3.050 0.390 ;
        RECT  1.240 -0.165 2.860 0.165 ;
        RECT  1.050 -0.165 1.240 0.300 ;
        RECT  0.220 -0.165 1.050 0.165 ;
        RECT  0.075 -0.165 0.220 0.545 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.005 1.110 4.125 1.965 ;
        RECT  3.370 1.635 4.005 1.965 ;
        RECT  3.370 1.390 3.650 1.490 ;
        RECT  3.230 1.390 3.370 1.965 ;
        RECT  2.940 1.390 3.230 1.490 ;
        RECT  0.770 1.635 3.230 1.965 ;
        RECT  0.770 1.390 1.020 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.310 1.390 0.630 1.485 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 0.510 3.895 0.675 ;
        RECT  3.750 1.110 3.895 1.290 ;
        RECT  3.195 0.510 3.250 0.675 ;
        RECT  3.195 1.110 3.250 1.290 ;
        RECT  2.950 0.785 3.235 0.885 ;
        RECT  2.850 0.500 2.950 1.300 ;
        RECT  2.750 0.500 2.850 0.590 ;
        RECT  1.350 1.210 2.850 1.300 ;
        RECT  1.235 1.390 2.830 1.490 ;
        RECT  2.660 0.310 2.750 0.590 ;
        RECT  1.540 0.310 2.660 0.410 ;
        RECT  1.450 0.310 1.540 0.480 ;
        RECT  0.520 0.390 1.450 0.480 ;
        RECT  1.135 1.210 1.235 1.490 ;
        RECT  0.195 1.210 1.135 1.300 ;
        RECT  0.075 1.210 0.195 1.450 ;
    END
END AO32D4

MACRO AO33D0
    CLASS CORE ;
    FOREIGN AO33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.275 2.150 1.490 ;
        RECT  2.015 0.275 2.050 0.480 ;
        RECT  2.015 1.255 2.050 1.490 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.910 1.950 1.090 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.090 ;
        RECT  0.990 0.700 1.050 0.950 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 0.700 0.830 0.950 ;
        RECT  0.650 0.700 0.760 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 -0.165 2.200 0.165 ;
        RECT  1.650 -0.165 1.840 0.410 ;
        RECT  0.235 -0.165 1.650 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.830 1.635 2.200 1.965 ;
        RECT  1.695 1.250 1.830 1.965 ;
        RECT  0.000 1.635 1.695 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.790 0.500 1.900 0.750 ;
        RECT  1.015 0.500 1.790 0.590 ;
        RECT  1.415 1.210 1.550 1.450 ;
        RECT  1.020 1.210 1.415 1.300 ;
        RECT  0.910 1.210 1.020 1.525 ;
        RECT  0.875 0.275 1.015 0.590 ;
        RECT  0.305 1.435 0.910 1.525 ;
        RECT  0.350 0.500 0.875 0.590 ;
        RECT  0.350 1.210 0.795 1.345 ;
        RECT  0.260 0.500 0.350 1.345 ;
        RECT  0.185 1.210 0.260 1.345 ;
        RECT  0.075 1.210 0.185 1.490 ;
    END
END AO33D0

MACRO AO33D1
    CLASS CORE ;
    FOREIGN AO33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.015 0.275 2.150 1.490 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.600 0.950 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.815 -0.165 2.200 0.165 ;
        RECT  1.625 -0.165 1.815 0.410 ;
        RECT  0.235 -0.165 1.625 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.635 2.200 1.965 ;
        RECT  1.680 1.100 1.810 1.965 ;
        RECT  1.265 1.635 1.680 1.965 ;
        RECT  1.075 1.390 1.265 1.965 ;
        RECT  0.000 1.635 1.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.800 0.500 1.900 0.950 ;
        RECT  0.350 0.500 1.800 0.590 ;
        RECT  0.960 1.210 1.535 1.300 ;
        RECT  0.860 1.210 0.960 1.490 ;
        RECT  0.295 1.390 0.860 1.490 ;
        RECT  0.350 1.210 0.745 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 1.210 0.260 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO33D1

MACRO AO33D2
    CLASS CORE ;
    FOREIGN AO33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.535 2.150 1.195 ;
        RECT  2.050 0.275 2.060 1.490 ;
        RECT  1.960 0.275 2.050 0.675 ;
        RECT  1.960 1.045 2.050 1.490 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.600 0.950 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.165 2.400 0.165 ;
        RECT  2.210 -0.165 2.330 0.455 ;
        RECT  1.790 -0.165 2.210 0.165 ;
        RECT  1.600 -0.165 1.790 0.410 ;
        RECT  0.235 -0.165 1.600 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.635 2.400 1.965 ;
        RECT  2.210 1.325 2.330 1.965 ;
        RECT  1.780 1.635 2.210 1.965 ;
        RECT  1.660 1.100 1.780 1.965 ;
        RECT  1.265 1.635 1.660 1.965 ;
        RECT  1.075 1.390 1.265 1.965 ;
        RECT  0.000 1.635 1.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.750 0.500 1.850 0.950 ;
        RECT  0.350 0.500 1.750 0.590 ;
        RECT  0.960 1.210 1.535 1.300 ;
        RECT  0.860 1.210 0.960 1.490 ;
        RECT  0.295 1.390 0.860 1.490 ;
        RECT  0.350 1.210 0.750 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 1.210 0.260 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO33D2

MACRO AO33D4
    CLASS CORE ;
    FOREIGN AO33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.310 4.305 0.690 ;
        RECT  4.250 1.110 4.305 1.490 ;
        RECT  3.950 0.310 4.250 1.490 ;
        RECT  3.650 0.310 3.950 0.690 ;
        RECT  3.650 1.110 3.950 1.490 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.1101 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.500 1.580 1.100 ;
        RECT  0.180 0.500 1.450 0.590 ;
        RECT  0.050 0.500 0.180 1.100 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.700 1.350 1.100 ;
        RECT  0.560 1.010 1.240 1.100 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.700 1.150 0.900 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.500 3.160 1.100 ;
        RECT  1.950 0.500 3.050 0.590 ;
        RECT  1.830 0.500 1.950 0.920 ;
        RECT  1.775 0.700 1.830 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.820 0.700 2.950 1.100 ;
        RECT  2.150 1.010 2.820 1.100 ;
        RECT  2.040 0.700 2.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.700 2.550 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 -0.165 4.600 0.165 ;
        RECT  4.415 -0.165 4.535 0.690 ;
        RECT  0.245 -0.165 4.415 0.165 ;
        RECT  0.055 -0.165 0.245 0.390 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 1.635 4.600 1.965 ;
        RECT  4.415 1.110 4.535 1.965 ;
        RECT  0.485 1.635 4.415 1.965 ;
        RECT  0.295 1.390 0.485 1.965 ;
        RECT  0.000 1.635 0.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 0.310 3.850 0.690 ;
        RECT  3.650 1.110 3.850 1.490 ;
        RECT  3.425 0.800 3.760 0.900 ;
        RECT  3.305 0.310 3.425 1.300 ;
        RECT  1.700 1.390 3.315 1.490 ;
        RECT  0.830 0.310 3.305 0.410 ;
        RECT  1.815 1.210 3.305 1.300 ;
        RECT  1.600 1.210 1.700 1.490 ;
        RECT  0.180 1.210 1.600 1.300 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END AO33D4

MACRO AOI211D0
    CLASS CORE ;
    FOREIGN AOI211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.090 ;
        RECT  0.980 0.500 1.250 0.590 ;
        RECT  0.865 0.280 0.980 0.590 ;
        RECT  0.355 0.500 0.865 0.590 ;
        RECT  0.355 1.215 0.485 1.325 ;
        RECT  0.265 0.500 0.355 1.325 ;
        RECT  0.195 0.500 0.265 0.590 ;
        RECT  0.065 0.310 0.195 0.590 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.155 1.090 ;
        RECT  0.970 0.700 1.045 0.950 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.760 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.165 1.400 0.165 ;
        RECT  1.150 -0.165 1.300 0.390 ;
        RECT  0.755 -0.165 1.150 0.165 ;
        RECT  0.555 -0.165 0.755 0.410 ;
        RECT  0.000 -0.165 0.555 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.635 1.400 1.965 ;
        RECT  1.150 1.245 1.300 1.965 ;
        RECT  0.000 1.635 1.150 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 1.240 0.715 1.525 ;
        RECT  0.175 1.435 0.605 1.525 ;
        RECT  0.065 1.240 0.175 1.525 ;
    END
END AOI211D0

MACRO AOI211D1
    CLASS CORE ;
    FOREIGN AOI211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.300 ;
        RECT  0.045 0.500 1.250 0.590 ;
        RECT  0.305 1.210 1.250 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.970 0.700 1.050 0.950 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.165 1.400 0.165 ;
        RECT  1.150 -0.165 1.300 0.390 ;
        RECT  0.755 -0.165 1.150 0.165 ;
        RECT  0.555 -0.165 0.755 0.410 ;
        RECT  0.000 -0.165 0.555 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.635 1.400 1.965 ;
        RECT  1.150 1.410 1.300 1.965 ;
        RECT  0.000 1.635 1.150 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.190 1.390 0.755 1.490 ;
        RECT  0.070 1.240 0.190 1.490 ;
    END
END AOI211D1

MACRO AOI211D2
    CLASS CORE ;
    FOREIGN AOI211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4420 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.500 2.355 1.290 ;
        RECT  0.300 0.500 2.245 0.600 ;
        RECT  1.340 1.200 2.245 1.290 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.710 1.150 1.090 ;
        RECT  0.170 1.000 1.030 1.090 ;
        RECT  0.050 0.700 0.170 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.710 2.150 1.090 ;
        RECT  1.370 1.000 2.045 1.090 ;
        RECT  1.250 0.710 1.370 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.955 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.165 2.400 0.165 ;
        RECT  0.770 0.310 1.280 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.045 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.635 2.400 1.965 ;
        RECT  0.560 1.390 0.750 1.965 ;
        RECT  0.000 1.635 0.560 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 1.400 2.310 1.505 ;
        RECT  1.125 1.210 1.225 1.505 ;
        RECT  0.185 1.210 1.125 1.300 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AOI211D2

MACRO AOI211D4
    CLASS CORE ;
    FOREIGN AOI211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9670 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.500 4.460 0.610 ;
        RECT  1.450 1.210 2.350 1.300 ;
        RECT  1.150 0.500 1.450 1.300 ;
        RECT  0.340 0.500 1.150 0.610 ;
        RECT  0.070 1.210 1.150 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.775 0.710 4.550 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 3.395 0.890 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2197 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 2.395 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 1.030 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 -0.165 4.800 0.165 ;
        RECT  3.570 0.300 4.730 0.410 ;
        RECT  3.430 -0.165 3.570 0.410 ;
        RECT  0.000 -0.165 3.430 0.165 ;
        RECT  2.460 0.300 3.430 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.175 1.635 4.800 1.965 ;
        RECT  4.175 1.390 4.470 1.490 ;
        RECT  4.035 1.390 4.175 1.965 ;
        RECT  3.740 1.390 4.035 1.490 ;
        RECT  0.000 1.635 4.035 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.550 0.500 4.460 0.610 ;
        RECT  1.550 1.210 2.350 1.300 ;
        RECT  0.340 0.500 1.050 0.610 ;
        RECT  0.070 1.210 1.050 1.300 ;
        RECT  2.460 1.210 4.720 1.300 ;
        RECT  0.330 1.390 3.430 1.490 ;
        RECT  0.225 0.300 2.370 0.410 ;
        RECT  0.105 0.300 0.225 0.560 ;
    END
END AOI211D4

MACRO AOI211XD0
    CLASS CORE ;
    FOREIGN AOI211XD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.090 ;
        RECT  0.980 0.500 1.250 0.590 ;
        RECT  0.870 0.280 0.980 0.590 ;
        RECT  0.355 0.500 0.870 0.590 ;
        RECT  0.355 1.215 0.495 1.325 ;
        RECT  0.265 0.500 0.355 1.325 ;
        RECT  0.195 0.500 0.265 0.590 ;
        RECT  0.070 0.310 0.195 0.590 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0434 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.155 1.090 ;
        RECT  0.970 0.700 1.045 0.950 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.760 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.165 1.400 0.165 ;
        RECT  1.150 -0.165 1.300 0.390 ;
        RECT  0.755 -0.165 1.150 0.165 ;
        RECT  0.555 -0.165 0.755 0.410 ;
        RECT  0.000 -0.165 0.555 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.635 1.400 1.965 ;
        RECT  1.150 1.245 1.300 1.965 ;
        RECT  0.000 1.635 1.150 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 1.240 0.715 1.525 ;
        RECT  0.175 1.435 0.605 1.525 ;
        RECT  0.065 1.240 0.175 1.525 ;
    END
END AOI211XD0

MACRO AOI211XD1
    CLASS CORE ;
    FOREIGN AOI211XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.510 2.350 1.300 ;
        RECT  0.855 0.510 2.240 0.600 ;
        RECT  1.375 1.200 2.240 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0861 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0860 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.090 ;
        RECT  0.355 1.000 1.045 1.090 ;
        RECT  0.245 0.710 0.355 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0860 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.550 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 -0.165 2.400 0.165 ;
        RECT  0.970 0.295 1.575 0.420 ;
        RECT  0.830 -0.165 0.970 0.420 ;
        RECT  0.000 -0.165 0.830 0.165 ;
        RECT  0.580 0.295 0.830 0.420 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.185 1.410 2.345 1.510 ;
        RECT  0.295 1.200 1.065 1.300 ;
        RECT  0.075 1.200 0.185 1.510 ;
    END
END AOI211XD1

MACRO AOI211XD2
    CLASS CORE ;
    FOREIGN AOI211XD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.500 3.845 0.600 ;
        RECT  1.155 1.110 2.045 1.290 ;
        RECT  1.045 0.500 1.155 1.290 ;
        RECT  0.795 0.500 1.045 0.600 ;
        RECT  0.295 1.110 1.045 1.290 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1726 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.710 3.950 0.925 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1716 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.925 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1724 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.925 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1716 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.370 -0.165 4.600 0.165 ;
        RECT  3.370 0.295 4.105 0.410 ;
        RECT  3.230 -0.165 3.370 0.410 ;
        RECT  0.000 -0.165 3.230 0.165 ;
        RECT  2.615 0.295 3.230 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.410 1.000 4.520 1.490 ;
        RECT  4.020 1.200 4.410 1.300 ;
        RECT  3.910 1.035 4.020 1.490 ;
        RECT  3.520 1.200 3.910 1.300 ;
        RECT  3.410 1.000 3.520 1.300 ;
        RECT  2.375 1.200 3.410 1.300 ;
        RECT  2.265 1.390 3.345 1.490 ;
        RECT  2.155 1.000 2.265 1.490 ;
        RECT  0.185 1.390 2.155 1.490 ;
        RECT  0.545 0.310 1.795 0.410 ;
        RECT  0.075 1.000 0.185 1.490 ;
    END
END AOI211XD2

MACRO AOI211XD4
    CLASS CORE ;
    FOREIGN AOI211XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.3000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 7.460 0.610 ;
        RECT  2.250 1.200 4.125 1.300 ;
        RECT  1.950 0.510 2.250 1.300 ;
        RECT  1.325 0.510 1.950 0.610 ;
        RECT  0.295 1.200 1.950 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.3432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.840 0.710 8.370 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.3432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.710 6.180 0.890 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.3449 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 3.980 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 1.765 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.680 -0.165 8.800 0.165 ;
        RECT  7.570 -0.165 7.680 0.585 ;
        RECT  6.570 -0.165 7.570 0.165 ;
        RECT  6.570 0.315 7.215 0.415 ;
        RECT  6.430 -0.165 6.570 0.415 ;
        RECT  0.000 -0.165 6.430 0.165 ;
        RECT  5.225 0.315 6.430 0.415 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.500 1.635 8.800 1.965 ;
        RECT  8.310 1.390 8.500 1.965 ;
        RECT  7.980 1.635 8.310 1.965 ;
        RECT  7.790 1.390 7.980 1.965 ;
        RECT  7.460 1.635 7.790 1.965 ;
        RECT  7.270 1.390 7.460 1.965 ;
        RECT  6.940 1.635 7.270 1.965 ;
        RECT  6.750 1.390 6.940 1.965 ;
        RECT  0.000 1.635 6.750 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.510 7.460 0.610 ;
        RECT  2.350 1.200 4.125 1.300 ;
        RECT  1.325 0.510 1.850 0.610 ;
        RECT  0.295 1.200 1.850 1.300 ;
        RECT  8.610 1.000 8.720 1.490 ;
        RECT  8.200 1.200 8.610 1.300 ;
        RECT  8.090 1.000 8.200 1.490 ;
        RECT  7.680 1.200 8.090 1.300 ;
        RECT  7.570 1.035 7.680 1.490 ;
        RECT  7.160 1.200 7.570 1.300 ;
        RECT  7.050 1.000 7.160 1.490 ;
        RECT  6.640 1.200 7.050 1.300 ;
        RECT  6.530 1.000 6.640 1.300 ;
        RECT  4.455 1.200 6.530 1.300 ;
        RECT  4.345 1.390 6.465 1.490 ;
        RECT  4.235 1.000 4.345 1.490 ;
        RECT  0.185 1.390 4.235 1.490 ;
        RECT  1.055 0.315 3.355 0.415 ;
        RECT  0.075 1.000 0.185 1.490 ;
    END
END AOI211XD4

MACRO AOI21D0
    CLASS CORE ;
    FOREIGN AOI21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0940 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.460 1.150 1.090 ;
        RECT  0.750 0.460 1.050 0.560 ;
        RECT  0.590 0.275 0.750 0.560 ;
        RECT  0.355 0.460 0.590 0.560 ;
        RECT  0.355 1.215 0.485 1.325 ;
        RECT  0.265 0.460 0.355 1.325 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.680 0.810 0.950 ;
        RECT  0.645 0.680 0.755 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.680 0.555 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 -0.165 1.200 0.165 ;
        RECT  0.870 -0.165 1.020 0.370 ;
        RECT  0.175 -0.165 0.870 0.165 ;
        RECT  0.065 -0.165 0.175 0.475 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 1.635 1.200 1.965 ;
        RECT  0.885 1.240 1.005 1.965 ;
        RECT  0.000 1.635 0.885 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 1.240 0.715 1.525 ;
        RECT  0.175 1.435 0.605 1.525 ;
        RECT  0.065 1.240 0.175 1.525 ;
    END
END AOI21D0

MACRO AOI21D1
    CLASS CORE ;
    FOREIGN AOI21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.460 1.150 1.300 ;
        RECT  0.565 0.460 1.050 0.560 ;
        RECT  0.305 1.210 1.050 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.810 0.950 ;
        RECT  0.650 0.680 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.165 1.200 0.165 ;
        RECT  0.860 -0.165 1.030 0.350 ;
        RECT  0.190 -0.165 0.860 0.165 ;
        RECT  0.070 -0.165 0.190 0.475 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.635 1.200 1.965 ;
        RECT  0.870 1.410 1.020 1.965 ;
        RECT  0.000 1.635 0.870 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.190 1.390 0.755 1.490 ;
        RECT  0.070 1.240 0.190 1.490 ;
    END
END AOI21D1

MACRO AOI21D2
    CLASS CORE ;
    FOREIGN AOI21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4100 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.565 0.500 1.755 0.590 ;
        RECT  0.565 1.210 1.505 1.300 ;
        RECT  0.450 0.500 0.565 1.300 ;
        RECT  0.045 0.500 0.450 0.590 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.700 0.360 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.350 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  0.950 1.010 1.450 1.100 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.750 0.700 0.850 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.245 -0.165 1.800 0.165 ;
        RECT  1.055 -0.165 1.245 0.410 ;
        RECT  0.000 -0.165 1.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.615 1.250 1.735 1.490 ;
        RECT  0.185 1.390 1.615 1.490 ;
        RECT  0.065 1.250 0.185 1.490 ;
    END
END AOI21D2

MACRO AOI21D4
    CLASS CORE ;
    FOREIGN AOI21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8010 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.500 0.500 3.305 0.600 ;
        RECT  2.400 0.500 2.500 1.300 ;
        RECT  0.850 1.210 2.400 1.300 ;
        RECT  0.850 0.500 1.030 0.590 ;
        RECT  0.550 0.500 0.850 1.300 ;
        RECT  0.320 0.500 0.550 0.590 ;
        RECT  0.050 1.210 0.550 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.770 3.370 0.900 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2197 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.770 2.240 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.355 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 -0.165 3.600 0.165 ;
        RECT  3.415 -0.165 3.535 0.675 ;
        RECT  2.535 -0.165 3.415 0.165 ;
        RECT  2.345 -0.165 2.535 0.410 ;
        RECT  0.000 -0.165 2.345 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 1.635 3.600 1.965 ;
        RECT  3.415 1.115 3.535 1.965 ;
        RECT  0.000 1.635 3.415 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.500 0.500 3.305 0.600 ;
        RECT  2.400 0.500 2.500 1.300 ;
        RECT  0.950 1.210 2.400 1.300 ;
        RECT  0.950 0.500 1.030 0.590 ;
        RECT  0.320 0.500 0.450 0.590 ;
        RECT  0.050 1.210 0.450 1.300 ;
        RECT  3.150 1.010 3.270 1.490 ;
        RECT  2.755 1.390 3.150 1.490 ;
        RECT  2.645 1.010 2.755 1.490 ;
        RECT  0.320 1.390 2.645 1.490 ;
        RECT  1.245 0.500 2.275 0.600 ;
        RECT  1.145 0.310 1.245 0.600 ;
        RECT  0.205 0.310 1.145 0.410 ;
        RECT  0.085 0.310 0.205 0.560 ;
    END
END AOI21D4

MACRO AOI221D0
    CLASS CORE ;
    FOREIGN AOI221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.310 1.445 0.425 ;
        RECT  0.950 1.090 1.075 1.220 ;
        RECT  0.850 1.090 0.950 1.305 ;
        RECT  0.350 1.215 0.850 1.305 ;
        RECT  0.350 0.310 0.550 0.490 ;
        RECT  0.250 0.310 0.350 1.305 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.160 1.090 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0285 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.530 1.550 1.235 ;
        RECT  0.760 0.530 1.440 0.620 ;
        RECT  0.660 0.530 0.760 0.700 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.600 0.550 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0291 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.960 0.930 ;
        RECT  0.755 0.820 0.850 0.930 ;
        RECT  0.650 0.820 0.755 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.710 1.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 1.345 1.520 1.515 ;
        RECT  0.270 1.410 1.390 1.515 ;
    END
END AOI221D0

MACRO AOI221D1
    CLASS CORE ;
    FOREIGN AOI221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 0.500 1.505 0.590 ;
        RECT  0.160 1.200 0.490 1.290 ;
        RECT  0.050 0.500 0.160 1.290 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 1.100 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.700 1.155 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.360 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.755 0.930 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.360 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.735 0.590 ;
        RECT  0.995 -0.165 1.615 0.165 ;
        RECT  0.820 -0.165 0.995 0.410 ;
        RECT  0.000 -0.165 0.820 0.165 ;
        RECT  0.550 0.295 0.820 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 1.635 1.800 1.965 ;
        RECT  1.615 1.210 1.735 1.965 ;
        RECT  0.000 1.635 1.615 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.795 1.390 1.505 1.500 ;
        RECT  0.705 1.210 1.245 1.300 ;
        RECT  0.605 1.110 0.705 1.500 ;
        RECT  0.050 1.400 0.605 1.500 ;
    END
END AOI221D1

MACRO AOI221D2
    CLASS CORE ;
    FOREIGN AOI221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.500 3.150 1.300 ;
        RECT  0.045 0.500 3.050 0.590 ;
        RECT  1.900 1.210 3.050 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.700 0.360 1.100 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.350 0.900 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.750 1.100 ;
        RECT  0.950 1.010 1.650 1.100 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.765 0.700 0.850 0.920 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.700 2.750 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.700 2.950 1.100 ;
        RECT  2.150 1.010 2.850 1.100 ;
        RECT  2.040 0.700 2.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.165 3.200 0.165 ;
        RECT  2.420 -0.165 2.610 0.410 ;
        RECT  0.770 -0.165 2.420 0.165 ;
        RECT  0.770 0.310 1.280 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.290 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.635 3.200 1.965 ;
        RECT  0.300 1.390 0.490 1.965 ;
        RECT  0.000 1.635 0.300 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.810 1.390 2.880 1.490 ;
        RECT  0.185 1.210 1.790 1.300 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AOI221D2

MACRO AOI221D4
    CLASS CORE ;
    FOREIGN AOI221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.515 2.640 0.685 ;
        RECT  2.250 1.110 2.595 1.490 ;
        RECT  1.950 0.515 2.250 1.490 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.600 0.950 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.700 0.950 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.355 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.570 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 -0.165 3.200 0.165 ;
        RECT  0.850 -0.165 1.000 0.410 ;
        RECT  0.245 -0.165 0.850 0.165 ;
        RECT  0.055 -0.165 0.245 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.635 3.200 1.965 ;
        RECT  2.750 1.335 2.860 1.965 ;
        RECT  1.815 1.635 2.750 1.965 ;
        RECT  1.680 1.110 1.815 1.965 ;
        RECT  0.000 1.635 1.680 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.515 2.640 0.685 ;
        RECT  2.350 1.110 2.595 1.490 ;
        RECT  3.115 0.310 3.155 1.210 ;
        RECT  3.045 0.310 3.115 1.490 ;
        RECT  2.965 0.310 3.045 0.410 ;
        RECT  3.015 1.110 3.045 1.490 ;
        RECT  2.775 1.110 3.015 1.210 ;
        RECT  2.865 0.500 2.955 0.945 ;
        RECT  2.855 0.500 2.865 0.590 ;
        RECT  2.755 0.295 2.855 0.590 ;
        RECT  2.685 0.800 2.775 1.210 ;
        RECT  1.515 0.295 2.755 0.405 ;
        RECT  2.495 0.800 2.685 0.900 ;
        RECT  0.835 1.390 1.555 1.490 ;
        RECT  1.385 0.295 1.515 0.590 ;
        RECT  0.360 0.500 1.385 0.590 ;
        RECT  0.725 1.210 1.295 1.300 ;
        RECT  0.605 1.210 0.725 1.510 ;
        RECT  0.180 1.410 0.605 1.510 ;
        RECT  0.360 1.210 0.495 1.300 ;
        RECT  0.270 0.500 0.360 1.300 ;
        RECT  0.060 1.240 0.180 1.510 ;
    END
END AOI221D4

MACRO AOI221XD4
    CLASS CORE ;
    FOREIGN AOI221XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.615 1.015 5.725 1.490 ;
        RECT  4.755 1.015 5.615 1.125 ;
        RECT  4.755 0.500 5.505 0.610 ;
        RECT  4.645 0.500 4.755 1.125 ;
        RECT  3.250 1.015 4.645 1.125 ;
        RECT  2.950 0.500 3.250 1.125 ;
        RECT  1.245 0.500 2.950 0.610 ;
        RECT  1.055 0.500 1.245 0.700 ;
        RECT  0.185 0.500 1.055 0.610 ;
        RECT  0.075 0.310 0.185 0.610 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2192 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.925 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.925 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.750 0.925 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.710 4.350 0.925 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.165 5.800 0.165 ;
        RECT  0.295 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 1.635 5.800 1.965 ;
        RECT  0.815 1.395 1.005 1.965 ;
        RECT  0.485 1.635 0.815 1.965 ;
        RECT  0.295 1.395 0.485 1.965 ;
        RECT  0.000 1.635 0.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.615 1.015 5.725 1.490 ;
        RECT  4.755 1.015 5.615 1.125 ;
        RECT  4.755 0.500 5.505 0.610 ;
        RECT  4.645 0.500 4.755 1.125 ;
        RECT  3.350 1.015 4.645 1.125 ;
        RECT  1.245 0.500 2.850 0.610 ;
        RECT  1.055 0.500 1.245 0.700 ;
        RECT  0.185 0.500 1.055 0.610 ;
        RECT  0.075 0.310 0.185 0.610 ;
        RECT  5.615 0.310 5.725 0.610 ;
        RECT  3.680 0.310 5.615 0.410 ;
        RECT  1.405 1.395 5.505 1.485 ;
        RECT  3.580 0.310 3.680 0.700 ;
        RECT  1.260 0.310 3.490 0.410 ;
        RECT  1.265 1.215 3.425 1.305 ;
        RECT  1.155 1.000 1.265 1.490 ;
        RECT  0.705 1.215 1.155 1.305 ;
        RECT  0.595 1.035 0.705 1.490 ;
        RECT  0.185 1.215 0.595 1.305 ;
        RECT  0.075 1.000 0.185 1.490 ;
    END
END AOI221XD4

MACRO AOI222D0
    CLASS CORE ;
    FOREIGN AOI222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1310 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.355 0.310 1.745 0.420 ;
        RECT  1.350 1.070 1.460 1.200 ;
        RECT  1.250 1.070 1.350 1.305 ;
        RECT  0.355 1.215 1.250 1.305 ;
        RECT  0.250 0.310 0.355 1.305 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.675 0.160 1.090 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.560 1.090 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0285 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.530 1.950 1.235 ;
        RECT  1.135 0.530 1.840 0.620 ;
        RECT  0.965 0.530 1.135 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.765 0.800 0.950 0.930 ;
        RECT  0.755 0.800 0.765 1.090 ;
        RECT  0.650 0.710 0.755 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.710 1.360 0.915 ;
        RECT  1.155 0.780 1.225 0.915 ;
        RECT  1.050 0.780 1.155 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.710 1.750 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.790 1.345 1.920 1.525 ;
        RECT  0.060 1.415 1.790 1.525 ;
    END
END AOI222D0

MACRO AOI222D1
    CLASS CORE ;
    FOREIGN AOI222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.510 1.585 0.600 ;
        RECT  0.150 1.200 0.515 1.290 ;
        RECT  0.050 0.510 0.150 1.290 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.700 1.950 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.160 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.950 1.100 ;
        RECT  0.790 0.710 0.850 0.950 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.710 0.605 0.950 ;
        RECT  0.450 0.710 0.550 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.035 -0.165 2.200 0.165 ;
        RECT  1.915 -0.165 2.035 0.590 ;
        RECT  0.770 -0.165 1.915 0.165 ;
        RECT  0.770 0.300 1.305 0.400 ;
        RECT  0.630 -0.165 0.770 0.400 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.065 0.300 0.630 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.635 2.200 1.965 ;
        RECT  1.770 1.390 2.095 1.500 ;
        RECT  1.630 1.390 1.770 1.965 ;
        RECT  1.395 1.390 1.630 1.500 ;
        RECT  0.000 1.635 1.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.845 1.210 1.835 1.300 ;
        RECT  0.065 1.400 1.285 1.510 ;
    END
END AOI222D1

MACRO AOI222D2
    CLASS CORE ;
    FOREIGN AOI222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5550 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.500 3.555 1.300 ;
        RECT  0.525 0.500 3.450 0.590 ;
        RECT  2.495 1.210 3.450 1.300 ;
        RECT  2.375 1.060 2.495 1.300 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.700 1.050 0.920 ;
        RECT  0.850 0.700 0.960 1.100 ;
        RECT  0.170 1.010 0.850 1.100 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.700 2.150 1.100 ;
        RECT  1.350 1.010 2.050 1.100 ;
        RECT  1.250 0.700 1.350 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.900 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.700 3.150 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.700 3.350 1.100 ;
        RECT  2.750 1.010 3.250 1.100 ;
        RECT  2.635 0.710 2.750 1.100 ;
        RECT  2.540 0.710 2.635 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.570 -0.165 3.600 0.165 ;
        RECT  2.570 0.310 3.060 0.410 ;
        RECT  2.430 -0.165 2.570 0.410 ;
        RECT  0.770 -0.165 2.430 0.165 ;
        RECT  2.065 0.310 2.430 0.410 ;
        RECT  0.770 0.310 1.235 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.045 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 1.390 3.305 1.490 ;
        RECT  0.185 1.210 2.265 1.300 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AOI222D2

MACRO AOI222D4
    CLASS CORE ;
    FOREIGN AOI222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.510 2.840 0.690 ;
        RECT  2.450 1.110 2.795 1.490 ;
        RECT  2.150 0.510 2.450 1.490 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.700 1.950 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.155 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.775 0.700 0.850 0.950 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.165 3.400 0.165 ;
        RECT  0.770 0.310 1.280 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.060 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.635 3.400 1.965 ;
        RECT  2.935 1.335 3.080 1.965 ;
        RECT  2.040 1.635 2.935 1.965 ;
        RECT  1.930 1.335 2.040 1.965 ;
        RECT  1.380 1.390 1.930 1.490 ;
        RECT  0.000 1.635 1.930 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.510 2.840 0.690 ;
        RECT  2.550 1.110 2.795 1.490 ;
        RECT  3.315 0.310 3.355 1.210 ;
        RECT  3.245 0.310 3.315 1.490 ;
        RECT  3.165 0.310 3.245 0.410 ;
        RECT  3.215 1.110 3.245 1.490 ;
        RECT  2.975 1.110 3.215 1.210 ;
        RECT  3.065 0.500 3.155 0.945 ;
        RECT  3.055 0.500 3.065 0.590 ;
        RECT  2.955 0.310 3.055 0.590 ;
        RECT  2.885 0.800 2.975 1.210 ;
        RECT  1.535 0.310 2.955 0.400 ;
        RECT  2.695 0.800 2.885 0.900 ;
        RECT  0.820 1.210 1.820 1.300 ;
        RECT  1.400 0.310 1.535 0.590 ;
        RECT  0.360 0.500 1.400 0.590 ;
        RECT  0.060 1.390 1.270 1.490 ;
        RECT  0.360 1.210 0.510 1.300 ;
        RECT  0.260 0.500 0.360 1.300 ;
    END
END AOI222D4

MACRO AOI222XD4
    CLASS CORE ;
    FOREIGN AOI222XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.815 1.015 6.925 1.490 ;
        RECT  4.450 1.015 6.815 1.125 ;
        RECT  4.450 0.500 6.705 0.610 ;
        RECT  4.150 0.500 4.450 1.125 ;
        RECT  1.295 0.500 4.150 0.610 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.395 0.710 0.805 0.890 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.395 0.710 1.805 0.890 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.710 3.005 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.595 0.710 4.005 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.195 0.710 5.605 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.195 0.710 6.605 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 7.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.045 1.635 7.000 1.965 ;
        RECT  1.855 1.395 2.045 1.965 ;
        RECT  1.525 1.635 1.855 1.965 ;
        RECT  1.335 1.395 1.525 1.965 ;
        RECT  1.005 1.635 1.335 1.965 ;
        RECT  0.815 1.395 1.005 1.965 ;
        RECT  0.485 1.635 0.815 1.965 ;
        RECT  0.295 1.395 0.485 1.965 ;
        RECT  0.000 1.635 0.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.815 1.015 6.925 1.490 ;
        RECT  4.550 1.015 6.815 1.125 ;
        RECT  4.550 0.500 6.705 0.610 ;
        RECT  1.295 0.500 4.050 0.610 ;
        RECT  6.815 0.300 6.925 0.610 ;
        RECT  4.705 0.300 6.815 0.410 ;
        RECT  2.615 1.395 6.705 1.485 ;
        RECT  2.505 1.215 4.625 1.305 ;
        RECT  2.365 0.300 4.615 0.410 ;
        RECT  2.395 1.020 2.505 1.490 ;
        RECT  2.265 1.215 2.395 1.305 ;
        RECT  2.155 1.020 2.265 1.490 ;
        RECT  1.185 0.300 2.255 0.410 ;
        RECT  1.745 1.215 2.155 1.305 ;
        RECT  1.635 1.035 1.745 1.490 ;
        RECT  1.225 1.215 1.635 1.305 ;
        RECT  1.115 1.000 1.225 1.490 ;
        RECT  1.075 0.275 1.185 0.670 ;
        RECT  0.705 1.215 1.115 1.305 ;
        RECT  0.185 0.300 1.075 0.410 ;
        RECT  0.595 1.035 0.705 1.490 ;
        RECT  0.185 1.215 0.595 1.305 ;
        RECT  0.075 0.275 0.185 0.670 ;
        RECT  0.075 1.000 0.185 1.490 ;
    END
END AOI222XD4

MACRO AOI22D0
    CLASS CORE ;
    FOREIGN AOI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.255 0.450 1.350 1.300 ;
        RECT  1.240 0.280 1.255 1.300 ;
        RECT  1.050 0.280 1.240 0.560 ;
        RECT  1.020 1.210 1.240 1.300 ;
        RECT  0.210 0.450 1.050 0.560 ;
        RECT  0.830 1.210 1.020 1.345 ;
        RECT  0.050 0.275 0.210 0.560 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.680 0.555 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.680 0.800 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.680 1.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 -0.165 1.400 0.165 ;
        RECT  0.580 -0.165 0.750 0.345 ;
        RECT  0.000 -0.165 0.580 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.715 1.435 1.335 1.525 ;
        RECT  0.615 1.210 0.715 1.525 ;
        RECT  0.210 1.210 0.615 1.300 ;
        RECT  0.080 1.210 0.210 1.450 ;
    END
END AOI22D0

MACRO AOI22D1
    CLASS CORE ;
    FOREIGN AOI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.460 1.350 1.290 ;
        RECT  0.050 0.460 1.240 0.560 ;
        RECT  0.830 1.200 1.240 1.290 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.680 0.550 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.680 0.810 0.950 ;
        RECT  0.650 0.680 0.750 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.680 1.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 -0.165 1.400 0.165 ;
        RECT  0.580 -0.165 0.750 0.345 ;
        RECT  0.000 -0.165 0.580 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 1.635 1.400 1.965 ;
        RECT  0.310 1.390 0.500 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.715 1.400 1.290 1.500 ;
        RECT  0.615 1.210 0.715 1.500 ;
        RECT  0.195 1.210 0.615 1.300 ;
        RECT  0.075 1.210 0.195 1.450 ;
    END
END AOI22D1

MACRO AOI22D2
    CLASS CORE ;
    FOREIGN AOI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.500 2.350 1.290 ;
        RECT  0.560 0.500 2.240 0.590 ;
        RECT  1.340 1.200 2.240 1.290 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.700 1.150 1.100 ;
        RECT  0.170 1.010 1.030 1.100 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.700 2.150 1.090 ;
        RECT  1.370 1.000 2.040 1.090 ;
        RECT  1.250 0.700 1.370 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.950 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.165 2.400 0.165 ;
        RECT  0.770 0.310 1.280 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.050 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.635 2.400 1.965 ;
        RECT  0.770 1.390 1.010 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.300 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 1.400 2.320 1.500 ;
        RECT  1.125 1.210 1.225 1.500 ;
        RECT  0.185 1.210 1.125 1.300 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AOI22D2

MACRO AOI22D4
    CLASS CORE ;
    FOREIGN AOI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.500 4.505 0.590 ;
        RECT  3.795 0.500 3.955 1.120 ;
        RECT  2.150 1.030 3.795 1.120 ;
        RECT  2.050 1.030 2.150 1.300 ;
        RECT  0.850 1.210 2.050 1.300 ;
        RECT  0.850 0.500 1.005 0.590 ;
        RECT  0.550 0.500 0.850 1.300 ;
        RECT  0.295 0.500 0.550 0.590 ;
        RECT  0.045 1.210 0.550 1.300 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.710 3.350 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.710 4.570 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.710 2.150 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.355 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.735 1.635 4.800 1.965 ;
        RECT  4.615 1.095 4.735 1.965 ;
        RECT  3.970 1.635 4.615 1.965 ;
        RECT  3.970 1.390 4.255 1.490 ;
        RECT  3.830 1.390 3.970 1.965 ;
        RECT  3.525 1.390 3.830 1.490 ;
        RECT  2.970 1.635 3.830 1.965 ;
        RECT  2.970 1.390 3.215 1.490 ;
        RECT  2.830 1.390 2.970 1.965 ;
        RECT  2.495 1.390 2.830 1.490 ;
        RECT  0.000 1.635 2.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.955 0.500 4.505 0.590 ;
        RECT  3.795 0.500 3.955 1.120 ;
        RECT  2.150 1.030 3.795 1.120 ;
        RECT  2.050 1.030 2.150 1.300 ;
        RECT  0.950 1.210 2.050 1.300 ;
        RECT  0.950 0.500 1.005 0.590 ;
        RECT  0.295 0.500 0.450 0.590 ;
        RECT  0.045 1.210 0.450 1.300 ;
        RECT  4.615 0.310 4.735 0.560 ;
        RECT  3.245 0.310 4.615 0.410 ;
        RECT  2.385 1.210 4.505 1.300 ;
        RECT  3.055 0.310 3.245 0.610 ;
        RECT  2.745 0.310 3.055 0.410 ;
        RECT  2.555 0.310 2.745 0.610 ;
        RECT  2.285 1.210 2.385 1.490 ;
        RECT  0.295 1.390 2.285 1.490 ;
        RECT  2.055 0.310 2.245 0.610 ;
        RECT  1.745 0.310 2.055 0.410 ;
        RECT  1.555 0.310 1.745 0.610 ;
        RECT  0.180 0.310 1.555 0.410 ;
        RECT  0.060 0.310 0.180 0.560 ;
    END
END AOI22D4

MACRO AOI31D0
    CLASS CORE ;
    FOREIGN AOI31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1480 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.510 1.350 1.100 ;
        RECT  0.965 0.510 1.240 0.600 ;
        RECT  0.810 0.285 0.965 0.600 ;
        RECT  0.350 0.510 0.810 0.600 ;
        RECT  0.640 1.075 0.750 1.375 ;
        RECT  0.350 1.275 0.640 1.375 ;
        RECT  0.260 0.510 0.350 1.375 ;
        RECT  0.190 1.275 0.260 1.375 ;
        RECT  0.050 1.275 0.190 1.490 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.150 1.100 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.550 1.165 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.930 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 -0.165 1.400 0.165 ;
        RECT  1.090 -0.165 1.265 0.400 ;
        RECT  0.235 -0.165 1.090 0.165 ;
        RECT  0.055 -0.165 0.235 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.635 1.400 1.965 ;
        RECT  1.140 1.255 1.280 1.965 ;
        RECT  0.000 1.635 1.140 1.965 ;
        END
    END VDD
END AOI31D0

MACRO AOI31D1
    CLASS CORE ;
    FOREIGN AOI31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2650 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.300 ;
        RECT  0.785 0.500 1.250 0.590 ;
        RECT  0.045 1.210 1.250 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 -0.165 1.400 0.165 ;
        RECT  1.090 -0.165 1.260 0.390 ;
        RECT  0.205 -0.165 1.090 0.165 ;
        RECT  0.075 -0.165 0.205 0.565 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.635 1.400 1.965 ;
        RECT  1.110 1.410 1.280 1.965 ;
        RECT  0.000 1.635 1.110 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.285 1.390 1.000 1.490 ;
    END
END AOI31D1

MACRO AOI31D2
    CLASS CORE ;
    FOREIGN AOI31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.390 2.350 1.100 ;
        RECT  1.350 0.390 2.250 0.480 ;
        RECT  1.550 1.010 2.250 1.100 ;
        RECT  1.450 1.010 1.550 1.300 ;
        RECT  0.310 1.210 1.450 1.300 ;
        RECT  1.250 0.310 1.350 0.480 ;
        RECT  0.790 0.310 1.250 0.410 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.900 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.780 1.665 0.890 ;
        RECT  1.450 0.570 1.550 0.890 ;
        RECT  1.150 0.570 1.450 0.660 ;
        RECT  1.050 0.500 1.150 0.660 ;
        RECT  0.360 0.500 1.050 0.590 ;
        RECT  0.270 0.500 0.360 0.780 ;
        RECT  0.170 0.680 0.270 0.780 ;
        RECT  0.050 0.680 0.170 1.120 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.775 1.350 1.100 ;
        RECT  0.550 1.010 1.250 1.100 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.700 0.950 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.785 -0.165 2.400 0.165 ;
        RECT  1.595 -0.165 1.785 0.300 ;
        RECT  0.180 -0.165 1.595 0.165 ;
        RECT  0.060 -0.165 0.180 0.570 ;
        RECT  0.000 -0.165 0.060 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.060 1.635 2.400 1.965 ;
        RECT  1.870 1.390 2.060 1.965 ;
        RECT  0.000 1.635 1.870 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.175 1.210 2.295 1.450 ;
        RECT  1.755 1.210 2.175 1.300 ;
        RECT  1.655 1.210 1.755 1.490 ;
        RECT  0.195 1.390 1.655 1.490 ;
        RECT  0.075 1.240 0.195 1.490 ;
    END
END AOI31D2

MACRO AOI31D4
    CLASS CORE ;
    FOREIGN AOI31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9870 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.555 0.500 4.290 0.590 ;
        RECT  3.445 0.500 3.555 1.150 ;
        RECT  3.150 1.040 3.445 1.150 ;
        RECT  3.050 1.040 3.150 1.300 ;
        RECT  1.050 1.210 3.050 1.300 ;
        RECT  0.750 0.500 1.050 1.300 ;
        RECT  0.295 0.500 0.750 0.590 ;
        RECT  0.045 1.210 0.750 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2206 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.775 4.355 0.900 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 3.200 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.710 2.020 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.710 0.630 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 -0.165 4.600 0.165 ;
        RECT  4.400 -0.165 4.520 0.685 ;
        RECT  0.000 -0.165 4.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.555 0.500 4.290 0.590 ;
        RECT  3.445 0.500 3.555 1.150 ;
        RECT  3.150 1.040 3.445 1.150 ;
        RECT  3.050 1.040 3.150 1.300 ;
        RECT  1.150 1.210 3.050 1.300 ;
        RECT  0.295 0.500 0.650 0.590 ;
        RECT  0.045 1.210 0.650 1.300 ;
        RECT  4.410 1.010 4.530 1.490 ;
        RECT  4.020 1.390 4.410 1.490 ;
        RECT  3.910 1.010 4.020 1.490 ;
        RECT  0.295 1.390 3.910 1.490 ;
        RECT  1.335 0.500 3.290 0.590 ;
        RECT  0.185 0.310 2.305 0.410 ;
        RECT  0.065 0.310 0.185 0.560 ;
    END
END AOI31D4

MACRO AOI32D0
    CLASS CORE ;
    FOREIGN AOI32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 0.280 0.965 0.600 ;
        RECT  0.150 0.510 0.825 0.600 ;
        RECT  0.180 1.210 0.795 1.345 ;
        RECT  0.150 1.210 0.180 1.490 ;
        RECT  0.050 0.510 0.150 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.700 1.395 0.950 ;
        RECT  1.250 0.700 1.350 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.150 1.095 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.350 1.095 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.580 1.095 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.950 1.095 ;
        RECT  0.740 0.710 0.850 0.950 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.165 1.600 0.165 ;
        RECT  1.370 -0.165 1.500 0.465 ;
        RECT  0.250 -0.165 1.370 0.165 ;
        RECT  0.065 -0.165 0.250 0.400 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.395 1.210 1.525 1.450 ;
        RECT  1.015 1.210 1.395 1.300 ;
        RECT  0.905 1.210 1.015 1.525 ;
        RECT  0.300 1.435 0.905 1.525 ;
    END
END AOI32D0

MACRO AOI32D1
    CLASS CORE ;
    FOREIGN AOI32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.310 0.960 0.600 ;
        RECT  0.150 0.510 0.835 0.600 ;
        RECT  0.150 1.210 0.750 1.300 ;
        RECT  0.050 0.510 0.150 1.300 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.700 1.395 0.950 ;
        RECT  1.250 0.700 1.350 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.150 1.100 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.350 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.580 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.950 1.100 ;
        RECT  0.740 0.710 0.850 0.950 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 -0.165 1.600 0.165 ;
        RECT  1.365 -0.165 1.505 0.585 ;
        RECT  0.250 -0.165 1.365 0.165 ;
        RECT  0.065 -0.165 0.250 0.400 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.635 1.600 1.965 ;
        RECT  1.080 1.390 1.270 1.965 ;
        RECT  0.000 1.635 1.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.385 1.210 1.505 1.450 ;
        RECT  0.965 1.210 1.385 1.300 ;
        RECT  0.865 1.210 0.965 1.500 ;
        RECT  0.290 1.390 0.865 1.500 ;
    END
END AOI32D1

MACRO AOI32D2
    CLASS CORE ;
    FOREIGN AOI32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.300 2.950 1.300 ;
        RECT  1.540 0.300 2.850 0.410 ;
        RECT  1.350 1.210 2.850 1.300 ;
        RECT  1.450 0.300 1.540 0.480 ;
        RECT  0.520 0.390 1.450 0.480 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.700 1.065 0.920 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.170 1.010 0.850 1.100 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.775 2.625 0.945 ;
        RECT  2.445 0.510 2.555 1.100 ;
        RECT  1.750 0.510 2.445 0.600 ;
        RECT  1.660 0.510 1.750 0.660 ;
        RECT  1.350 0.570 1.660 0.660 ;
        RECT  1.235 0.570 1.350 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.355 1.100 ;
        RECT  1.575 1.010 2.250 1.100 ;
        RECT  1.450 0.775 1.575 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 -0.165 3.000 0.165 ;
        RECT  1.050 -0.165 1.240 0.300 ;
        RECT  0.215 -0.165 1.050 0.165 ;
        RECT  0.075 -0.165 0.215 0.545 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.635 3.000 1.965 ;
        RECT  0.770 1.390 1.025 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.310 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.235 1.390 2.840 1.490 ;
        RECT  1.135 1.210 1.235 1.490 ;
        RECT  0.200 1.210 1.135 1.300 ;
        RECT  0.080 1.210 0.200 1.450 ;
    END
END AOI32D2

MACRO AOI32D4
    CLASS CORE ;
    FOREIGN AOI32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.510 2.900 0.675 ;
        RECT  2.650 1.110 2.900 1.290 ;
        RECT  2.350 0.510 2.650 1.290 ;
        RECT  2.200 0.510 2.350 0.675 ;
        RECT  2.200 1.110 2.350 1.290 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.700 1.395 0.950 ;
        RECT  1.250 0.700 1.350 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.700 1.150 1.100 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.580 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.740 0.700 0.850 0.950 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 -0.165 3.200 0.165 ;
        RECT  3.010 -0.165 3.130 0.675 ;
        RECT  2.370 -0.165 3.010 0.165 ;
        RECT  2.370 0.310 2.660 0.410 ;
        RECT  2.230 -0.165 2.370 0.410 ;
        RECT  1.530 -0.165 2.230 0.165 ;
        RECT  1.930 0.310 2.230 0.410 ;
        RECT  1.340 -0.165 1.530 0.410 ;
        RECT  0.240 -0.165 1.340 0.165 ;
        RECT  0.050 -0.165 0.240 0.410 ;
        RECT  0.000 -0.165 0.050 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.635 3.200 1.965 ;
        RECT  3.010 1.035 3.130 1.965 ;
        RECT  2.370 1.635 3.010 1.965 ;
        RECT  2.370 1.390 2.660 1.490 ;
        RECT  2.230 1.390 2.370 1.965 ;
        RECT  1.935 1.390 2.230 1.490 ;
        RECT  1.270 1.635 2.230 1.965 ;
        RECT  1.080 1.390 1.270 1.965 ;
        RECT  0.000 1.635 1.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 0.510 2.900 0.675 ;
        RECT  2.750 1.110 2.900 1.290 ;
        RECT  2.200 0.510 2.250 0.675 ;
        RECT  2.200 1.110 2.250 1.290 ;
        RECT  2.050 0.785 2.230 0.895 ;
        RECT  1.950 0.535 2.050 1.185 ;
        RECT  1.820 0.535 1.950 0.675 ;
        RECT  1.820 1.035 1.950 1.185 ;
        RECT  1.610 0.785 1.840 0.895 ;
        RECT  1.720 0.275 1.820 0.675 ;
        RECT  1.720 1.035 1.820 1.465 ;
        RECT  1.510 0.500 1.610 0.895 ;
        RECT  0.965 1.210 1.530 1.300 ;
        RECT  0.360 0.500 1.510 0.590 ;
        RECT  0.865 1.210 0.965 1.490 ;
        RECT  0.300 1.390 0.865 1.490 ;
        RECT  0.360 1.210 0.750 1.300 ;
        RECT  0.260 0.500 0.360 1.300 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AOI32D4

MACRO AOI32XD4
    CLASS CORE ;
    FOREIGN AOI32XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.1480 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.795 1.015 5.905 1.490 ;
        RECT  2.450 1.015 5.795 1.125 ;
        RECT  2.450 0.500 3.350 0.610 ;
        RECT  2.150 0.500 2.450 1.125 ;
        RECT  1.335 0.500 2.150 0.610 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.395 0.710 0.805 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.395 0.710 1.805 0.890 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.995 0.710 5.405 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.795 0.710 4.205 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.795 0.710 3.205 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.370 -0.165 6.000 0.165 ;
        RECT  5.370 0.300 5.700 0.410 ;
        RECT  5.230 -0.165 5.370 0.410 ;
        RECT  0.770 -0.165 5.230 0.165 ;
        RECT  4.975 0.300 5.230 0.410 ;
        RECT  0.770 0.300 1.005 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.295 0.300 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.305 1.635 6.000 1.965 ;
        RECT  2.115 1.395 2.305 1.965 ;
        RECT  1.785 1.635 2.115 1.965 ;
        RECT  1.595 1.395 1.785 1.965 ;
        RECT  1.265 1.635 1.595 1.965 ;
        RECT  1.075 1.395 1.265 1.965 ;
        RECT  0.745 1.635 1.075 1.965 ;
        RECT  0.555 1.395 0.745 1.965 ;
        RECT  0.185 1.635 0.555 1.965 ;
        RECT  0.075 1.035 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.795 1.015 5.905 1.490 ;
        RECT  2.550 1.015 5.795 1.125 ;
        RECT  2.550 0.500 3.350 0.610 ;
        RECT  1.335 0.500 2.050 0.610 ;
        RECT  3.650 0.500 5.935 0.610 ;
        RECT  2.005 1.215 5.685 1.305 ;
        RECT  2.385 0.300 4.645 0.410 ;
        RECT  1.225 0.300 2.295 0.410 ;
        RECT  1.895 1.035 2.005 1.490 ;
        RECT  1.485 1.215 1.895 1.305 ;
        RECT  1.375 1.035 1.485 1.490 ;
        RECT  0.965 1.215 1.375 1.305 ;
        RECT  1.115 0.275 1.225 0.670 ;
        RECT  0.185 0.500 1.115 0.610 ;
        RECT  0.855 1.035 0.965 1.490 ;
        RECT  0.445 1.215 0.855 1.305 ;
        RECT  0.335 1.035 0.445 1.490 ;
        RECT  0.075 0.275 0.185 0.670 ;
    END
END AOI32XD4

MACRO AOI33D0
    CLASS CORE ;
    FOREIGN AOI33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1410 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.310 0.985 0.490 ;
        RECT  0.565 1.200 0.745 1.345 ;
        RECT  0.350 1.200 0.565 1.290 ;
        RECT  0.260 0.310 0.350 1.290 ;
        RECT  0.250 0.310 0.260 0.490 ;
        RECT  0.185 1.200 0.260 1.290 ;
        RECT  0.050 1.200 0.185 1.490 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 1.090 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.700 1.150 1.090 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0289 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0285 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0285 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.700 0.800 0.950 ;
        RECT  0.645 0.700 0.755 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.165 1.800 0.165 ;
        RECT  1.600 -0.165 1.735 0.480 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.295 1.725 1.965 ;
        RECT  0.000 1.635 1.615 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.355 1.210 1.465 1.450 ;
        RECT  0.965 1.210 1.355 1.300 ;
        RECT  0.855 1.210 0.965 1.525 ;
        RECT  0.475 1.435 0.855 1.525 ;
        RECT  0.295 1.380 0.475 1.525 ;
    END
END AOI33D0

MACRO AOI33D1
    CLASS CORE ;
    FOREIGN AOI33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2650 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.310 0.985 0.490 ;
        RECT  0.350 1.210 0.745 1.300 ;
        RECT  0.260 0.310 0.350 1.300 ;
        RECT  0.250 0.310 0.260 0.490 ;
        RECT  0.045 1.210 0.260 1.300 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 1.100 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.700 1.150 1.100 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.800 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.735 0.570 ;
        RECT  0.000 -0.165 1.615 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 1.635 1.800 1.965 ;
        RECT  1.615 1.230 1.735 1.965 ;
        RECT  0.000 1.635 1.615 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.295 1.390 1.505 1.490 ;
    END
END AOI33D1

MACRO AOI33D2
    CLASS CORE ;
    FOREIGN AOI33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.310 3.350 1.190 ;
        RECT  2.880 0.310 3.250 0.400 ;
        RECT  3.070 1.100 3.250 1.190 ;
        RECT  2.980 1.100 3.070 1.300 ;
        RECT  1.850 1.210 2.980 1.300 ;
        RECT  0.825 0.310 2.880 0.405 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.500 1.580 1.100 ;
        RECT  0.350 0.500 1.450 0.590 ;
        RECT  0.205 0.500 0.350 1.100 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.700 1.350 1.100 ;
        RECT  0.560 1.010 1.240 1.100 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.700 1.150 0.900 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.035 0.510 3.150 0.990 ;
        RECT  1.950 0.510 3.035 0.600 ;
        RECT  1.815 0.510 1.950 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.750 0.710 2.865 0.930 ;
        RECT  2.650 0.710 2.750 1.100 ;
        RECT  2.160 1.010 2.650 1.100 ;
        RECT  2.050 0.710 2.160 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.550 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.260 -0.165 3.400 0.165 ;
        RECT  0.070 -0.165 0.260 0.410 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.635 3.400 1.965 ;
        RECT  0.770 1.390 1.035 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.310 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.190 1.300 3.300 1.490 ;
        RECT  1.735 1.390 3.190 1.490 ;
        RECT  1.635 1.210 1.735 1.490 ;
        RECT  0.195 1.210 1.635 1.300 ;
        RECT  0.075 1.210 0.195 1.450 ;
    END
END AOI33D2

MACRO AOI33D4
    CLASS CORE ;
    FOREIGN AOI33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.515 2.640 0.685 ;
        RECT  2.250 1.110 2.595 1.490 ;
        RECT  1.950 0.515 2.250 1.490 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.600 0.950 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.700 1.350 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.945 0.700 1.050 0.950 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.800 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.240 -0.165 3.200 0.165 ;
        RECT  0.050 -0.165 0.240 0.410 ;
        RECT  0.000 -0.165 0.050 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.635 3.200 1.965 ;
        RECT  2.750 1.335 2.860 1.965 ;
        RECT  1.805 1.635 2.750 1.965 ;
        RECT  1.695 1.000 1.805 1.965 ;
        RECT  1.080 1.390 1.695 1.490 ;
        RECT  0.000 1.635 1.695 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.515 2.640 0.685 ;
        RECT  2.350 1.110 2.595 1.490 ;
        RECT  3.115 0.310 3.155 1.210 ;
        RECT  3.045 0.310 3.115 1.490 ;
        RECT  2.965 0.310 3.045 0.410 ;
        RECT  3.015 1.110 3.045 1.490 ;
        RECT  2.775 1.110 3.015 1.210 ;
        RECT  2.865 0.500 2.955 0.945 ;
        RECT  2.855 0.500 2.865 0.590 ;
        RECT  2.755 0.295 2.855 0.590 ;
        RECT  2.685 0.795 2.775 1.210 ;
        RECT  0.490 0.295 2.755 0.405 ;
        RECT  2.445 0.795 2.685 0.905 ;
        RECT  0.965 1.210 1.530 1.300 ;
        RECT  0.865 1.210 0.965 1.490 ;
        RECT  0.300 1.390 0.865 1.490 ;
        RECT  0.350 1.210 0.750 1.300 ;
        RECT  0.380 0.295 0.490 0.590 ;
        RECT  0.350 0.500 0.380 0.590 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.065 1.210 0.185 1.450 ;
    END
END AOI33D4

MACRO AOI33XD4
    CLASS CORE ;
    FOREIGN AOI33XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.1150 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.015 1.015 7.125 1.490 ;
        RECT  3.850 1.015 7.015 1.125 ;
        RECT  3.850 0.500 4.605 0.610 ;
        RECT  3.550 0.500 3.850 1.125 ;
        RECT  2.595 0.500 3.550 0.610 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.395 0.710 0.805 0.890 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.595 0.710 2.005 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.710 3.005 0.890 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.210 0.710 6.605 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.995 0.710 5.405 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.995 0.710 4.405 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 7.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.565 1.635 7.200 1.965 ;
        RECT  3.375 1.395 3.565 1.965 ;
        RECT  3.045 1.635 3.375 1.965 ;
        RECT  2.855 1.395 3.045 1.965 ;
        RECT  2.525 1.635 2.855 1.965 ;
        RECT  2.335 1.395 2.525 1.965 ;
        RECT  2.005 1.635 2.335 1.965 ;
        RECT  1.815 1.395 2.005 1.965 ;
        RECT  1.370 1.635 1.815 1.965 ;
        RECT  1.370 1.395 1.505 1.505 ;
        RECT  1.230 1.395 1.370 1.965 ;
        RECT  1.065 1.395 1.230 1.505 ;
        RECT  0.745 1.635 1.230 1.965 ;
        RECT  0.555 1.395 0.745 1.965 ;
        RECT  0.185 1.635 0.555 1.965 ;
        RECT  0.075 1.035 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.015 1.015 7.125 1.490 ;
        RECT  3.950 1.015 7.015 1.125 ;
        RECT  3.950 0.500 4.605 0.610 ;
        RECT  2.595 0.500 3.450 0.610 ;
        RECT  7.015 0.275 7.125 0.670 ;
        RECT  6.125 0.500 7.015 0.610 ;
        RECT  3.265 1.215 6.905 1.305 ;
        RECT  6.015 0.275 6.125 0.670 ;
        RECT  4.935 0.500 6.015 0.610 ;
        RECT  4.825 0.300 5.905 0.410 ;
        RECT  4.715 0.275 4.825 0.670 ;
        RECT  3.645 0.300 4.715 0.410 ;
        RECT  2.485 0.300 3.555 0.410 ;
        RECT  3.155 1.035 3.265 1.490 ;
        RECT  2.745 1.215 3.155 1.305 ;
        RECT  2.635 1.035 2.745 1.490 ;
        RECT  2.225 1.215 2.635 1.305 ;
        RECT  2.375 0.275 2.485 0.670 ;
        RECT  1.295 0.300 2.375 0.410 ;
        RECT  1.185 0.500 2.265 0.610 ;
        RECT  2.115 1.035 2.225 1.490 ;
        RECT  1.705 1.215 2.115 1.305 ;
        RECT  1.595 1.035 1.705 1.490 ;
        RECT  0.965 1.215 1.595 1.305 ;
        RECT  1.075 0.275 1.185 0.670 ;
        RECT  0.185 0.500 1.075 0.610 ;
        RECT  0.855 1.035 0.965 1.490 ;
        RECT  0.445 1.215 0.855 1.305 ;
        RECT  0.335 1.035 0.445 1.490 ;
        RECT  0.075 0.275 0.185 0.670 ;
    END
END AOI33XD4

MACRO BENCD1
    CLASS CORE ;
    FOREIGN BENCD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.275 0.175 0.645 ;
        RECT  0.150 1.055 0.175 1.490 ;
        RECT  0.050 0.275 0.150 1.490 ;
        END
    END X2
    PIN S
        ANTENNADIFFAREA 0.2320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.510 4.090 0.600 ;
        RECT  3.550 1.025 3.750 1.115 ;
        RECT  3.440 0.510 3.550 1.115 ;
        END
    END S
    PIN M2
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.700 3.350 0.890 ;
        END
    END M2
    PIN M1
        ANTENNAGATEAREA 0.1408 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 0.710 2.550 0.890 ;
        RECT  2.040 0.510 2.150 0.890 ;
        RECT  1.855 0.510 2.040 0.600 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0870 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.710 1.950 0.890 ;
        RECT  1.550 0.710 1.640 0.945 ;
        RECT  1.195 0.855 1.550 0.945 ;
        END
    END M0
    PIN A
        ANTENNADIFFAREA 0.2000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.645 0.510 2.755 1.115 ;
        RECT  2.260 0.510 2.645 0.600 ;
        RECT  2.440 1.025 2.645 1.115 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.475 -0.165 4.400 0.165 ;
        RECT  3.305 -0.165 3.475 0.400 ;
        RECT  2.975 -0.165 3.305 0.165 ;
        RECT  2.845 -0.165 2.975 0.390 ;
        RECT  1.535 -0.165 2.845 0.165 ;
        RECT  1.405 -0.165 1.535 0.425 ;
        RECT  0.435 -0.165 1.405 0.165 ;
        RECT  0.335 -0.165 0.435 0.445 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.330 1.635 4.400 1.965 ;
        RECT  4.220 1.055 4.330 1.965 ;
        RECT  1.545 1.635 4.220 1.965 ;
        RECT  1.375 1.395 1.545 1.965 ;
        RECT  0.435 1.635 1.375 1.965 ;
        RECT  0.345 1.240 0.435 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.195 0.290 4.305 0.600 ;
        RECT  3.565 0.290 4.195 0.400 ;
        RECT  4.040 0.725 4.130 1.495 ;
        RECT  1.895 1.405 4.040 1.495 ;
        RECT  3.860 0.725 3.950 1.315 ;
        RECT  3.700 0.725 3.860 0.895 ;
        RECT  2.095 1.225 3.860 1.315 ;
        RECT  2.935 0.500 3.225 0.590 ;
        RECT  2.935 1.025 3.150 1.115 ;
        RECT  2.845 0.500 2.935 1.115 ;
        RECT  2.525 0.295 2.710 0.410 ;
        RECT  1.975 0.295 2.525 0.385 ;
        RECT  2.005 1.035 2.095 1.315 ;
        RECT  1.035 1.035 2.005 1.125 ;
        RECT  1.805 1.215 1.895 1.495 ;
        RECT  1.735 0.295 1.835 0.385 ;
        RECT  0.835 1.215 1.805 1.305 ;
        RECT  1.645 0.295 1.735 0.620 ;
        RECT  1.405 0.530 1.645 0.620 ;
        RECT  1.315 0.530 1.405 0.765 ;
        RECT  1.035 0.675 1.315 0.765 ;
        RECT  1.115 0.400 1.205 0.585 ;
        RECT  0.835 0.495 1.115 0.585 ;
        RECT  0.945 0.675 1.035 1.125 ;
        RECT  0.635 1.395 1.015 1.505 ;
        RECT  0.635 0.315 1.000 0.405 ;
        RECT  0.745 0.495 0.835 1.305 ;
        RECT  0.510 0.750 0.745 0.920 ;
        RECT  0.545 0.315 0.635 0.640 ;
        RECT  0.545 1.030 0.635 1.505 ;
        RECT  0.355 0.550 0.545 0.640 ;
        RECT  0.355 1.030 0.545 1.120 ;
        RECT  0.265 0.550 0.355 1.120 ;
        RECT  0.250 0.750 0.265 0.920 ;
    END
END BENCD1

MACRO BENCD2
    CLASS CORE ;
    FOREIGN BENCD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.275 0.430 0.645 ;
        RECT  0.350 1.055 0.430 1.490 ;
        RECT  0.330 0.275 0.350 1.490 ;
        RECT  0.250 0.510 0.330 1.310 ;
        END
    END X2
    PIN S
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.755 0.510 6.105 0.690 ;
        RECT  5.645 0.510 5.755 1.125 ;
        RECT  5.395 0.510 5.645 0.690 ;
        RECT  4.650 1.015 5.645 1.125 ;
        END
    END S
    PIN M2
        ANTENNAGATEAREA 0.1660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.895 ;
        END
    END M2
    PIN M1
        ANTENNAGATEAREA 0.1552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.710 3.150 0.890 ;
        RECT  2.350 0.710 2.840 0.800 ;
        RECT  2.250 0.510 2.350 0.800 ;
        RECT  2.065 0.510 2.250 0.600 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.1431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.160 0.925 ;
        RECT  1.425 0.835 1.850 0.925 ;
        END
    END M0
    PIN A
        ANTENNADIFFAREA 0.4150 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.555 1.035 4.085 1.125 ;
        RECT  3.445 0.510 3.555 1.125 ;
        RECT  2.460 0.510 3.445 0.600 ;
        RECT  3.415 1.035 3.445 1.125 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.040 -0.165 6.400 0.165 ;
        RECT  4.850 -0.165 5.040 0.480 ;
        RECT  4.210 -0.165 4.850 0.165 ;
        RECT  4.030 -0.165 4.210 0.415 ;
        RECT  1.775 -0.165 4.030 0.165 ;
        RECT  1.655 -0.165 1.775 0.425 ;
        RECT  0.000 -0.165 1.655 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.705 1.635 6.400 1.965 ;
        RECT  1.585 1.395 1.705 1.965 ;
        RECT  0.000 1.635 1.585 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.215 0.310 6.325 0.560 ;
        RECT  6.215 1.055 6.325 1.485 ;
        RECT  5.285 0.310 6.215 0.410 ;
        RECT  5.140 1.395 6.215 1.485 ;
        RECT  6.000 0.800 6.140 0.900 ;
        RECT  5.900 0.800 6.000 1.305 ;
        RECT  4.950 1.215 5.900 1.305 ;
        RECT  4.545 0.800 5.535 0.900 ;
        RECT  5.175 0.275 5.285 0.690 ;
        RECT  4.715 0.590 5.175 0.690 ;
        RECT  4.860 1.215 4.950 1.525 ;
        RECT  1.885 1.435 4.860 1.525 ;
        RECT  4.605 0.275 4.715 0.690 ;
        RECT  4.455 0.800 4.545 1.325 ;
        RECT  2.065 1.235 4.455 1.325 ;
        RECT  4.355 0.275 4.430 0.690 ;
        RECT  4.320 0.275 4.355 1.125 ;
        RECT  4.245 0.510 4.320 1.125 ;
        RECT  3.755 0.510 4.245 0.600 ;
        RECT  4.175 1.035 4.245 1.125 ;
        RECT  3.430 0.305 3.920 0.415 ;
        RECT  3.645 0.510 3.755 0.915 ;
        RECT  3.240 0.285 3.430 0.415 ;
        RECT  2.155 1.035 3.325 1.125 ;
        RECT  2.200 0.285 3.240 0.395 ;
        RECT  1.955 0.285 2.085 0.395 ;
        RECT  1.975 1.035 2.065 1.325 ;
        RECT  1.255 1.035 1.975 1.125 ;
        RECT  1.865 0.285 1.955 0.620 ;
        RECT  1.795 1.215 1.885 1.525 ;
        RECT  1.640 0.530 1.865 0.620 ;
        RECT  1.055 1.215 1.795 1.305 ;
        RECT  1.550 0.530 1.640 0.745 ;
        RECT  1.255 0.655 1.550 0.745 ;
        RECT  1.350 0.325 1.450 0.565 ;
        RECT  1.055 0.475 1.350 0.565 ;
        RECT  1.165 0.655 1.255 1.125 ;
        RECT  0.855 0.295 1.240 0.385 ;
        RECT  0.855 1.395 1.215 1.505 ;
        RECT  0.965 0.475 1.055 1.305 ;
        RECT  0.720 0.750 0.965 0.920 ;
        RECT  0.765 0.295 0.855 0.640 ;
        RECT  0.765 1.030 0.855 1.505 ;
        RECT  0.610 0.550 0.765 0.640 ;
        RECT  0.610 1.030 0.765 1.120 ;
        RECT  0.520 0.550 0.610 1.120 ;
        RECT  0.480 0.750 0.520 0.920 ;
    END
END BENCD2

MACRO BENCD4
    CLASS CORE ;
    FOREIGN BENCD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.310 0.940 0.690 ;
        RECT  0.650 1.110 0.940 1.490 ;
        RECT  0.350 0.310 0.650 1.490 ;
        RECT  0.295 0.310 0.350 0.690 ;
        RECT  0.295 1.110 0.350 1.490 ;
        END
    END X2
    PIN S
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.555 0.510 10.485 0.690 ;
        RECT  9.445 0.510 9.555 1.125 ;
        RECT  8.735 0.510 9.445 0.690 ;
        RECT  7.450 1.015 9.445 1.125 ;
        END
    END S
    PIN M2
        ANTENNAGATEAREA 0.3305 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.710 6.950 0.895 ;
        END
    END M2
    PIN M1
        ANTENNAGATEAREA 0.2595 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 0.710 5.195 0.890 ;
        RECT  3.365 0.710 4.400 0.800 ;
        RECT  3.275 0.510 3.365 0.800 ;
        RECT  3.060 0.510 3.275 0.600 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.2843 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 3.165 0.945 ;
        RECT  2.400 0.855 2.850 0.945 ;
        END
    END M0
    PIN A
        ANTENNADIFFAREA 0.7360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.755 1.035 6.705 1.125 ;
        RECT  5.645 0.510 5.755 1.125 ;
        RECT  3.455 0.510 5.645 0.600 ;
        RECT  5.515 1.035 5.645 1.125 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.385 -0.165 10.800 0.165 ;
        RECT  8.235 -0.165 8.385 0.500 ;
        RECT  7.865 -0.165 8.235 0.165 ;
        RECT  7.715 -0.165 7.865 0.500 ;
        RECT  7.295 -0.165 7.715 0.165 ;
        RECT  7.115 -0.165 7.295 0.415 ;
        RECT  6.785 -0.165 7.115 0.165 ;
        RECT  6.605 -0.165 6.785 0.415 ;
        RECT  2.785 -0.165 6.605 0.165 ;
        RECT  2.665 -0.165 2.785 0.425 ;
        RECT  2.265 -0.165 2.665 0.165 ;
        RECT  2.075 -0.165 2.265 0.385 ;
        RECT  0.185 -0.165 2.075 0.165 ;
        RECT  0.075 -0.165 0.185 0.690 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.930 1.635 10.800 1.965 ;
        RECT  7.740 1.395 7.930 1.965 ;
        RECT  2.760 1.635 7.740 1.965 ;
        RECT  2.650 1.405 2.760 1.965 ;
        RECT  2.210 1.635 2.650 1.965 ;
        RECT  2.060 1.405 2.210 1.965 ;
        RECT  0.185 1.635 2.060 1.965 ;
        RECT  0.075 1.110 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 0.310 0.940 0.690 ;
        RECT  0.750 1.110 0.940 1.490 ;
        RECT  10.585 1.055 10.715 1.485 ;
        RECT  10.595 0.310 10.705 0.560 ;
        RECT  8.625 0.310 10.595 0.410 ;
        RECT  10.205 1.395 10.585 1.485 ;
        RECT  9.750 0.800 10.500 0.900 ;
        RECT  10.055 1.055 10.205 1.485 ;
        RECT  8.475 1.395 10.055 1.485 ;
        RECT  9.650 0.800 9.750 1.305 ;
        RECT  7.600 1.215 9.650 1.305 ;
        RECT  7.345 0.800 9.100 0.900 ;
        RECT  8.515 0.275 8.625 0.690 ;
        RECT  8.105 0.590 8.515 0.690 ;
        RECT  7.995 0.275 8.105 0.690 ;
        RECT  7.585 0.590 7.995 0.690 ;
        RECT  7.500 1.215 7.600 1.525 ;
        RECT  7.475 0.275 7.585 0.690 ;
        RECT  2.940 1.435 7.500 1.525 ;
        RECT  7.255 0.800 7.345 1.325 ;
        RECT  3.120 1.235 7.255 1.325 ;
        RECT  7.060 0.510 7.165 1.125 ;
        RECT  6.350 0.510 7.060 0.600 ;
        RECT  6.970 1.035 7.060 1.125 ;
        RECT  5.935 0.305 6.495 0.415 ;
        RECT  6.250 0.510 6.350 0.860 ;
        RECT  5.910 0.760 6.250 0.860 ;
        RECT  5.845 0.305 5.935 0.650 ;
        RECT  5.465 0.305 5.845 0.415 ;
        RECT  5.275 0.285 5.465 0.415 ;
        RECT  3.215 1.035 5.425 1.125 ;
        RECT  3.205 0.285 5.275 0.395 ;
        RECT  3.030 1.035 3.120 1.325 ;
        RECT  2.965 0.285 3.085 0.395 ;
        RECT  2.905 1.035 3.030 1.135 ;
        RECT  2.875 0.285 2.965 0.620 ;
        RECT  2.850 1.225 2.940 1.525 ;
        RECT  2.060 1.035 2.905 1.125 ;
        RECT  2.740 0.530 2.875 0.620 ;
        RECT  2.525 1.225 2.850 1.315 ;
        RECT  2.650 0.530 2.740 0.765 ;
        RECT  2.060 0.675 2.650 0.765 ;
        RECT  1.960 0.495 2.540 0.585 ;
        RECT  2.335 1.215 2.525 1.315 ;
        RECT  1.565 1.215 2.335 1.305 ;
        RECT  1.930 0.675 2.060 1.125 ;
        RECT  1.860 0.325 1.960 0.585 ;
        RECT  1.565 0.495 1.860 0.585 ;
        RECT  1.140 0.295 1.750 0.385 ;
        RECT  1.140 1.395 1.705 1.505 ;
        RECT  1.475 0.495 1.565 1.305 ;
        RECT  1.250 0.745 1.475 0.915 ;
        RECT  1.050 0.295 1.140 1.505 ;
        RECT  0.855 0.800 1.050 0.910 ;
    END
END BENCD4

MACRO BHD
    CLASS CORE ;
    FOREIGN BHD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNAGATEAREA 0.0550 ;
        ANTENNADIFFAREA 0.0520 ;
        DIRECTION INOUT ;
        PORT
        LAYER M1 ;
        RECT  0.655 0.305 0.755 1.385 ;
        RECT  0.645 0.305 0.655 0.690 ;
        RECT  0.650 1.110 0.655 1.385 ;
        RECT  0.565 1.275 0.650 1.385 ;
        RECT  0.575 0.305 0.645 0.415 ;
        RECT  0.335 0.555 0.645 0.690 ;
        RECT  0.225 0.555 0.335 0.895 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 -0.165 0.800 0.165 ;
        RECT  0.335 -0.165 0.445 0.465 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 1.635 0.800 1.965 ;
        RECT  0.335 1.225 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.560 0.780 0.565 0.960 ;
        RECT  0.455 0.780 0.560 1.105 ;
        RECT  0.185 1.005 0.455 1.105 ;
        RECT  0.135 0.335 0.215 0.445 ;
        RECT  0.135 1.005 0.185 1.435 ;
        RECT  0.045 0.335 0.135 1.435 ;
    END
END BHD

MACRO BMLD1
    CLASS CORE ;
    FOREIGN BMLD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        ANTENNAGATEAREA 0.0944 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.215 0.710 4.350 1.095 ;
        END
    END X2
    PIN S
        ANTENNAGATEAREA 0.0523 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 0.890 ;
        RECT  1.550 0.710 1.650 0.890 ;
        END
    END S
    PIN PP
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.275 4.750 1.490 ;
        RECT  4.620 0.275 4.650 0.675 ;
        RECT  4.620 1.085 4.650 1.490 ;
        END
    END PP
    PIN M1
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.570 1.090 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0914 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.150 0.690 ;
        RECT  3.020 0.510 3.050 0.690 ;
        RECT  2.920 0.510 3.020 0.890 ;
        END
    END M0
    PIN A
        ANTENNAGATEAREA 0.0523 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.695 1.950 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.460 1.635 4.800 1.965 ;
        RECT  4.350 1.230 4.460 1.965 ;
        RECT  0.000 1.635 4.350 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.530 0.775 4.560 0.945 ;
        RECT  4.440 0.275 4.530 0.945 ;
        RECT  3.620 0.275 4.440 0.365 ;
        RECT  4.125 1.305 4.235 1.490 ;
        RECT  4.125 0.475 4.230 0.600 ;
        RECT  4.035 0.475 4.125 1.490 ;
        RECT  3.900 0.715 4.035 0.885 ;
        RECT  3.800 0.485 3.945 0.595 ;
        RECT  3.800 1.305 3.910 1.525 ;
        RECT  3.710 0.485 3.800 1.525 ;
        RECT  0.175 1.435 3.710 1.525 ;
        RECT  3.530 0.275 3.620 1.325 ;
        RECT  3.350 0.400 3.440 1.325 ;
        RECT  3.260 0.400 3.350 0.600 ;
        RECT  3.215 1.235 3.350 1.325 ;
        RECT  3.150 0.785 3.260 1.125 ;
        RECT  3.105 1.035 3.150 1.125 ;
        RECT  3.015 1.035 3.105 1.325 ;
        RECT  2.310 1.235 3.015 1.325 ;
        RECT  2.815 1.035 2.905 1.125 ;
        RECT  2.815 0.395 2.830 0.600 ;
        RECT  2.725 0.395 2.815 1.125 ;
        RECT  2.580 0.715 2.725 0.885 ;
        RECT  2.490 1.035 2.635 1.125 ;
        RECT  2.490 0.470 2.615 0.605 ;
        RECT  2.400 0.275 2.490 1.125 ;
        RECT  1.495 0.275 2.400 0.365 ;
        RECT  2.220 0.475 2.310 1.325 ;
        RECT  2.040 0.455 2.130 1.325 ;
        RECT  1.860 0.455 2.040 0.545 ;
        RECT  1.000 1.235 2.040 1.325 ;
        RECT  1.460 1.035 1.600 1.125 ;
        RECT  1.460 0.275 1.495 0.600 ;
        RECT  1.395 0.275 1.460 1.125 ;
        RECT  1.360 0.455 1.395 1.125 ;
        RECT  1.235 1.035 1.270 1.125 ;
        RECT  1.135 0.275 1.235 1.125 ;
        RECT  0.360 0.275 1.135 0.365 ;
        RECT  1.090 1.035 1.135 1.125 ;
        RECT  1.000 0.455 1.025 0.565 ;
        RECT  0.910 0.455 1.000 1.325 ;
        RECT  0.840 0.455 0.910 0.565 ;
        RECT  0.860 1.095 0.910 1.325 ;
        RECT  0.750 0.745 0.820 0.915 ;
        RECT  0.660 0.475 0.750 1.325 ;
        RECT  0.555 0.475 0.660 0.565 ;
        RECT  0.555 1.215 0.660 1.325 ;
        RECT  0.270 0.275 0.360 0.925 ;
        RECT  0.230 0.755 0.270 0.925 ;
        RECT  0.140 0.275 0.175 0.645 ;
        RECT  0.140 1.085 0.175 1.525 ;
        RECT  0.050 0.275 0.140 1.525 ;
    END
END BMLD1

MACRO BMLD2
    CLASS CORE ;
    FOREIGN BMLD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        ANTENNAGATEAREA 0.0947 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.215 0.710 4.350 1.095 ;
        END
    END X2
    PIN S
        ANTENNAGATEAREA 0.0523 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 0.890 ;
        RECT  1.550 0.710 1.650 0.890 ;
        END
    END S
    PIN PP
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.310 4.750 1.490 ;
        RECT  4.525 0.310 4.650 0.410 ;
        RECT  4.570 1.085 4.650 1.490 ;
        END
    END PP
    PIN M1
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.570 1.090 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0914 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.150 0.690 ;
        RECT  3.020 0.510 3.050 0.690 ;
        RECT  2.920 0.510 3.020 0.890 ;
        END
    END M0
    PIN A
        ANTENNAGATEAREA 0.0523 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.695 1.950 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.530 0.775 4.560 0.945 ;
        RECT  4.440 0.500 4.530 0.945 ;
        RECT  4.415 0.500 4.440 0.600 ;
        RECT  4.325 0.275 4.415 0.600 ;
        RECT  3.620 0.275 4.325 0.365 ;
        RECT  4.125 0.475 4.215 0.585 ;
        RECT  4.125 1.305 4.215 1.490 ;
        RECT  4.035 0.475 4.125 1.490 ;
        RECT  3.900 0.715 4.035 0.885 ;
        RECT  3.800 0.485 3.945 0.595 ;
        RECT  3.800 1.305 3.910 1.525 ;
        RECT  3.710 0.485 3.800 1.525 ;
        RECT  0.175 1.435 3.710 1.525 ;
        RECT  3.530 0.275 3.620 1.325 ;
        RECT  3.350 0.400 3.440 1.325 ;
        RECT  3.260 0.400 3.350 0.600 ;
        RECT  3.215 1.235 3.350 1.325 ;
        RECT  3.150 0.785 3.260 1.125 ;
        RECT  3.105 1.035 3.150 1.125 ;
        RECT  3.015 1.035 3.105 1.325 ;
        RECT  2.310 1.235 3.015 1.325 ;
        RECT  2.815 1.035 2.905 1.125 ;
        RECT  2.815 0.400 2.830 0.600 ;
        RECT  2.725 0.400 2.815 1.125 ;
        RECT  2.580 0.715 2.725 0.885 ;
        RECT  2.490 1.035 2.635 1.125 ;
        RECT  2.490 0.485 2.610 0.595 ;
        RECT  2.400 0.275 2.490 1.125 ;
        RECT  1.495 0.275 2.400 0.365 ;
        RECT  2.220 0.475 2.310 1.325 ;
        RECT  2.040 0.455 2.130 1.325 ;
        RECT  1.860 0.455 2.040 0.545 ;
        RECT  1.000 1.235 2.040 1.325 ;
        RECT  1.460 1.035 1.600 1.125 ;
        RECT  1.460 0.275 1.495 0.600 ;
        RECT  1.395 0.275 1.460 1.125 ;
        RECT  1.360 0.455 1.395 1.125 ;
        RECT  1.235 1.035 1.270 1.125 ;
        RECT  1.135 0.275 1.235 1.125 ;
        RECT  0.360 0.275 1.135 0.365 ;
        RECT  1.090 1.035 1.135 1.125 ;
        RECT  1.000 0.455 1.025 0.565 ;
        RECT  0.910 0.455 1.000 1.325 ;
        RECT  0.840 0.455 0.910 0.565 ;
        RECT  0.860 1.095 0.910 1.325 ;
        RECT  0.750 0.745 0.820 0.915 ;
        RECT  0.660 0.475 0.750 1.325 ;
        RECT  0.555 0.475 0.660 0.565 ;
        RECT  0.555 1.215 0.660 1.325 ;
        RECT  0.270 0.275 0.360 0.925 ;
        RECT  0.230 0.755 0.270 0.925 ;
        RECT  0.140 0.275 0.175 0.645 ;
        RECT  0.140 1.085 0.175 1.525 ;
        RECT  0.050 0.275 0.140 1.525 ;
    END
END BMLD2

MACRO BMLD4
    CLASS CORE ;
    FOREIGN BMLD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        ANTENNAGATEAREA 0.0938 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.765 6.150 1.290 ;
        RECT  5.880 0.765 6.050 0.955 ;
        END
    END X2
    PIN S
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.350 0.890 ;
        END
    END S
    PIN PP
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.310 6.900 0.690 ;
        RECT  6.850 1.110 6.900 1.490 ;
        RECT  6.550 0.310 6.850 1.490 ;
        RECT  6.210 0.310 6.550 0.490 ;
        RECT  6.260 1.110 6.550 1.490 ;
        END
    END PP
    PIN M1
        ANTENNAGATEAREA 0.0924 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 0.710 0.810 0.895 ;
        RECT  0.650 0.710 0.770 1.090 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0937 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.510 4.350 0.895 ;
        RECT  4.105 0.710 4.250 0.895 ;
        END
    END M0
    PIN A
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.750 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.120 -0.165 7.200 0.165 ;
        RECT  7.010 -0.165 7.120 0.690 ;
        RECT  0.180 -0.165 7.010 0.165 ;
        RECT  0.070 -0.165 0.180 0.645 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.125 1.635 7.200 1.965 ;
        RECT  7.015 1.110 7.125 1.965 ;
        RECT  6.140 1.635 7.015 1.965 ;
        RECT  5.950 1.390 6.140 1.965 ;
        RECT  0.180 1.635 5.950 1.965 ;
        RECT  0.070 1.085 0.180 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.210 0.310 6.450 0.490 ;
        RECT  6.260 1.110 6.450 1.490 ;
        RECT  6.260 0.585 6.360 0.945 ;
        RECT  6.080 0.585 6.260 0.675 ;
        RECT  5.990 0.275 6.080 0.675 ;
        RECT  5.285 0.275 5.990 0.365 ;
        RECT  5.790 0.485 5.880 0.595 ;
        RECT  5.790 1.110 5.840 1.490 ;
        RECT  5.700 0.485 5.790 1.490 ;
        RECT  5.565 0.725 5.700 0.895 ;
        RECT  5.465 0.485 5.610 0.595 ;
        RECT  5.465 1.305 5.580 1.525 ;
        RECT  5.375 0.485 5.465 1.525 ;
        RECT  0.435 1.435 5.375 1.525 ;
        RECT  5.195 0.275 5.285 1.325 ;
        RECT  5.015 0.385 5.105 1.325 ;
        RECT  4.555 0.385 5.015 0.515 ;
        RECT  4.405 1.235 5.015 1.325 ;
        RECT  4.445 0.310 4.555 0.515 ;
        RECT  4.450 0.710 4.550 1.125 ;
        RECT  4.295 1.035 4.450 1.125 ;
        RECT  4.205 1.035 4.295 1.325 ;
        RECT  3.500 1.235 4.205 1.325 ;
        RECT  4.005 1.035 4.095 1.125 ;
        RECT  3.980 0.465 4.080 0.575 ;
        RECT  3.980 0.810 4.005 1.125 ;
        RECT  3.915 0.465 3.980 1.125 ;
        RECT  3.890 0.465 3.915 0.895 ;
        RECT  3.770 0.725 3.890 0.895 ;
        RECT  3.680 1.035 3.825 1.125 ;
        RECT  3.680 0.470 3.800 0.595 ;
        RECT  3.590 0.275 3.680 1.125 ;
        RECT  2.230 0.275 3.590 0.365 ;
        RECT  3.410 0.475 3.500 1.325 ;
        RECT  3.230 0.455 3.320 1.325 ;
        RECT  2.540 0.455 3.230 0.545 ;
        RECT  1.240 1.235 3.230 1.325 ;
        RECT  1.745 1.035 2.325 1.125 ;
        RECT  2.090 0.275 2.230 0.550 ;
        RECT  1.745 0.275 2.090 0.365 ;
        RECT  1.625 0.275 1.745 1.125 ;
        RECT  1.375 0.275 1.510 1.125 ;
        RECT  0.685 0.275 1.375 0.365 ;
        RECT  1.330 1.035 1.375 1.125 ;
        RECT  1.240 0.455 1.265 0.565 ;
        RECT  1.150 0.455 1.240 1.325 ;
        RECT  1.080 0.455 1.150 0.565 ;
        RECT  1.100 1.095 1.150 1.325 ;
        RECT  0.990 0.745 1.060 0.915 ;
        RECT  0.900 0.475 0.990 1.325 ;
        RECT  0.795 0.475 0.900 0.565 ;
        RECT  0.795 1.215 0.900 1.325 ;
        RECT  0.595 0.275 0.685 0.600 ;
        RECT  0.560 0.500 0.595 0.600 ;
        RECT  0.470 0.500 0.560 0.935 ;
        RECT  0.380 0.310 0.485 0.410 ;
        RECT  0.380 1.085 0.435 1.525 ;
        RECT  0.290 0.310 0.380 1.525 ;
    END
END BMLD4

MACRO BUFFD0
    CLASS CORE ;
    FOREIGN BUFFD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 0.310 0.750 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.180 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 -0.165 0.800 0.165 ;
        RECT  0.315 -0.165 0.500 0.420 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.635 0.800 1.965 ;
        RECT  0.315 1.380 0.495 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.475 0.730 0.530 0.940 ;
        RECT  0.375 0.510 0.475 1.290 ;
        RECT  0.200 0.510 0.375 0.600 ;
        RECT  0.200 1.200 0.375 1.290 ;
        RECT  0.090 0.285 0.200 0.600 ;
        RECT  0.090 1.200 0.200 1.490 ;
    END
END BUFFD0

MACRO BUFFD1
    CLASS CORE ;
    FOREIGN BUFFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 0.310 0.750 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.180 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 -0.165 0.800 0.165 ;
        RECT  0.315 -0.165 0.500 0.420 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.635 0.800 1.965 ;
        RECT  0.315 1.380 0.495 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.475 0.730 0.530 0.940 ;
        RECT  0.375 0.510 0.475 1.290 ;
        RECT  0.200 0.510 0.375 0.600 ;
        RECT  0.200 1.200 0.375 1.290 ;
        RECT  0.090 0.280 0.200 0.600 ;
        RECT  0.090 1.200 0.200 1.490 ;
    END
END BUFFD1

MACRO BUFFD12
    CLASS CORE ;
    FOREIGN BUFFD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.0920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.325 4.105 0.690 ;
        RECT  2.850 1.100 4.105 1.475 ;
        RECT  2.350 0.325 2.850 1.475 ;
        RECT  1.335 0.325 2.350 0.690 ;
        RECT  1.335 1.100 2.350 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.355 0.710 0.815 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.705 ;
        RECT  0.185 -0.165 4.215 0.165 ;
        RECT  0.075 -0.165 0.185 0.705 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.095 4.325 1.965 ;
        RECT  0.185 1.635 4.215 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.325 4.105 0.690 ;
        RECT  2.950 1.100 4.105 1.475 ;
        RECT  1.335 0.325 2.250 0.690 ;
        RECT  1.335 1.100 2.250 1.475 ;
        RECT  3.010 0.800 4.140 0.940 ;
        RECT  1.225 0.800 2.190 0.940 ;
        RECT  1.075 0.470 1.225 1.190 ;
        RECT  0.995 0.470 1.075 0.620 ;
        RECT  0.975 1.040 1.075 1.190 ;
        RECT  0.825 0.285 0.995 0.620 ;
        RECT  0.845 1.040 0.975 1.500 ;
        RECT  0.455 1.040 0.845 1.190 ;
        RECT  0.475 0.470 0.825 0.620 ;
        RECT  0.305 0.285 0.475 0.620 ;
        RECT  0.325 1.040 0.455 1.500 ;
    END
END BUFFD12

MACRO BUFFD16
    CLASS CORE ;
    FOREIGN BUFFD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.4560 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.335 5.440 0.700 ;
        RECT  3.650 1.100 5.440 1.475 ;
        RECT  3.150 0.335 3.650 1.475 ;
        RECT  1.650 0.335 3.150 0.700 ;
        RECT  1.650 1.100 3.150 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2730 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.710 1.270 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 -0.165 5.800 0.165 ;
        RECT  5.550 -0.165 5.660 0.695 ;
        RECT  0.000 -0.165 5.550 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.635 5.800 1.965 ;
        RECT  5.550 1.040 5.660 1.965 ;
        RECT  0.000 1.635 5.550 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 0.335 5.440 0.700 ;
        RECT  3.750 1.100 5.440 1.475 ;
        RECT  1.650 0.335 3.050 0.700 ;
        RECT  1.650 1.100 3.050 1.475 ;
        RECT  3.915 0.810 5.505 0.950 ;
        RECT  1.540 0.810 2.915 0.950 ;
        RECT  1.360 0.400 1.540 1.340 ;
        RECT  0.080 0.400 1.360 0.580 ;
        RECT  0.080 1.160 1.360 1.340 ;
    END
END BUFFD16

MACRO BUFFD2
    CLASS CORE ;
    FOREIGN BUFFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.275 0.765 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.195 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.165 1.200 0.165 ;
        RECT  0.905 -0.165 1.015 0.695 ;
        RECT  0.500 -0.165 0.905 0.165 ;
        RECT  0.330 -0.165 0.500 0.390 ;
        RECT  0.000 -0.165 0.330 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 1.635 1.200 1.965 ;
        RECT  0.905 1.040 1.015 1.965 ;
        RECT  0.500 1.635 0.905 1.965 ;
        RECT  0.330 1.410 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.420 0.500 0.530 1.300 ;
        RECT  0.185 0.500 0.420 0.600 ;
        RECT  0.185 1.200 0.420 1.300 ;
        RECT  0.075 0.390 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.425 ;
    END
END BUFFD2

MACRO BUFFD20
    CLASS CORE ;
    FOREIGN BUFFD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.8200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.325 6.505 0.690 ;
        RECT  4.250 1.110 6.505 1.475 ;
        RECT  3.750 0.325 4.250 1.475 ;
        RECT  1.805 0.325 3.750 0.690 ;
        RECT  1.805 1.110 3.750 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3309 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.090 ;
        RECT  0.495 0.785 1.245 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 -0.165 6.800 0.165 ;
        RECT  6.615 -0.165 6.725 0.695 ;
        RECT  0.185 -0.165 6.615 0.165 ;
        RECT  0.075 -0.165 0.185 0.695 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 1.635 6.800 1.965 ;
        RECT  6.615 1.040 6.725 1.965 ;
        RECT  0.185 1.635 6.615 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.350 0.325 6.505 0.690 ;
        RECT  4.350 1.110 6.505 1.475 ;
        RECT  1.805 0.325 3.650 0.690 ;
        RECT  1.805 1.110 3.650 1.475 ;
        RECT  4.490 0.800 6.540 0.940 ;
        RECT  1.685 0.800 3.590 0.940 ;
        RECT  1.465 0.285 1.685 1.490 ;
        RECT  0.945 0.285 1.465 0.505 ;
        RECT  0.945 1.270 1.465 1.490 ;
        RECT  0.835 0.285 0.945 0.695 ;
        RECT  0.835 1.040 0.945 1.490 ;
        RECT  0.445 0.285 0.835 0.505 ;
        RECT  0.445 1.270 0.835 1.490 ;
        RECT  0.335 0.285 0.445 0.695 ;
        RECT  0.335 1.040 0.445 1.490 ;
    END
END BUFFD20

MACRO BUFFD24
    CLASS CORE ;
    FOREIGN BUFFD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 2.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.325 7.885 0.690 ;
        RECT  4.850 1.110 7.885 1.475 ;
        RECT  4.350 0.325 4.850 1.475 ;
        RECT  2.045 0.325 4.350 0.690 ;
        RECT  2.045 1.110 4.350 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3868 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 0.785 1.360 0.895 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.105 -0.165 8.200 0.165 ;
        RECT  7.995 -0.165 8.105 0.695 ;
        RECT  0.000 -0.165 7.995 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.105 1.635 8.200 1.965 ;
        RECT  7.995 1.020 8.105 1.965 ;
        RECT  0.000 1.635 7.995 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.950 0.325 7.885 0.690 ;
        RECT  4.950 1.110 7.885 1.475 ;
        RECT  2.045 0.325 4.250 0.690 ;
        RECT  2.045 1.110 4.250 1.475 ;
        RECT  5.135 0.800 7.875 0.940 ;
        RECT  1.730 0.800 4.190 0.940 ;
        RECT  1.480 0.285 1.730 1.505 ;
        RECT  1.190 0.285 1.480 0.535 ;
        RECT  1.190 1.255 1.480 1.505 ;
        RECT  1.070 0.285 1.190 0.685 ;
        RECT  1.070 1.040 1.190 1.505 ;
        RECT  0.690 0.285 1.070 0.535 ;
        RECT  0.690 1.255 1.070 1.505 ;
        RECT  0.570 0.285 0.690 0.685 ;
        RECT  0.570 1.040 0.690 1.505 ;
        RECT  0.075 0.285 0.570 0.535 ;
        RECT  0.075 1.255 0.570 1.505 ;
    END
END BUFFD24

MACRO BUFFD3
    CLASS CORE ;
    FOREIGN BUFFD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3270 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.275 1.350 1.490 ;
        RECT  0.805 0.650 1.215 0.950 ;
        RECT  0.695 0.275 0.805 1.470 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.355 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.065 -0.165 1.400 0.165 ;
        RECT  0.955 -0.165 1.065 0.540 ;
        RECT  0.585 -0.165 0.955 0.165 ;
        RECT  0.375 -0.165 0.585 0.410 ;
        RECT  0.000 -0.165 0.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.065 1.635 1.400 1.965 ;
        RECT  0.955 1.060 1.065 1.965 ;
        RECT  0.585 1.635 0.955 1.965 ;
        RECT  0.375 1.390 0.585 1.965 ;
        RECT  0.000 1.635 0.375 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.500 0.500 0.605 1.300 ;
        RECT  0.105 0.500 0.500 0.600 ;
        RECT  0.105 1.200 0.500 1.300 ;
    END
END BUFFD3

MACRO BUFFD4
    CLASS CORE ;
    FOREIGN BUFFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.345 0.275 1.455 1.470 ;
        RECT  1.150 0.505 1.345 1.210 ;
        RECT  0.955 0.505 1.150 0.675 ;
        RECT  0.955 1.040 1.150 1.210 ;
        RECT  0.840 0.275 0.955 0.675 ;
        RECT  0.845 1.040 0.955 1.470 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.785 0.505 0.890 ;
        RECT  0.050 0.700 0.155 1.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 -0.165 1.800 0.165 ;
        RECT  1.605 -0.165 1.715 0.695 ;
        RECT  0.195 -0.165 1.605 0.165 ;
        RECT  0.085 -0.165 0.195 0.525 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.635 1.800 1.965 ;
        RECT  1.605 1.020 1.715 1.965 ;
        RECT  0.195 1.635 1.605 1.965 ;
        RECT  0.085 1.260 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.505 1.050 0.675 ;
        RECT  0.955 1.040 1.050 1.210 ;
        RECT  0.840 0.275 0.955 0.675 ;
        RECT  0.845 1.040 0.955 1.470 ;
        RECT  0.730 0.785 0.925 0.890 ;
        RECT  0.630 0.585 0.730 1.150 ;
        RECT  0.455 0.585 0.630 0.695 ;
        RECT  0.455 1.040 0.630 1.150 ;
        RECT  0.345 0.275 0.455 0.695 ;
        RECT  0.345 1.040 0.455 1.470 ;
    END
END BUFFD4

MACRO BUFFD6
    CLASS CORE ;
    FOREIGN BUFFD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.5460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.310 2.075 0.690 ;
        RECT  1.650 1.110 2.075 1.490 ;
        RECT  1.350 0.310 1.650 1.490 ;
        RECT  0.845 0.310 1.350 0.690 ;
        RECT  0.845 1.110 1.350 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.785 0.525 0.890 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 -0.165 2.400 0.165 ;
        RECT  2.185 -0.165 2.295 0.695 ;
        RECT  0.735 -0.165 2.185 0.165 ;
        RECT  0.625 -0.165 0.735 0.475 ;
        RECT  0.215 -0.165 0.625 0.165 ;
        RECT  0.105 -0.165 0.215 0.475 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 1.635 2.400 1.965 ;
        RECT  2.185 1.020 2.295 1.965 ;
        RECT  0.735 1.635 2.185 1.965 ;
        RECT  0.625 1.260 0.735 1.965 ;
        RECT  0.215 1.635 0.625 1.965 ;
        RECT  0.105 1.260 0.215 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.750 0.310 2.075 0.690 ;
        RECT  1.750 1.110 2.075 1.490 ;
        RECT  0.845 0.310 1.250 0.690 ;
        RECT  0.845 1.110 1.250 1.490 ;
        RECT  0.735 0.785 1.225 0.890 ;
        RECT  0.635 0.585 0.735 1.150 ;
        RECT  0.475 0.585 0.635 0.695 ;
        RECT  0.475 1.040 0.635 1.150 ;
        RECT  0.365 0.275 0.475 0.695 ;
        RECT  0.365 1.040 0.475 1.470 ;
    END
END BUFFD6

MACRO BUFFD8
    CLASS CORE ;
    FOREIGN BUFFD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.325 2.850 0.690 ;
        RECT  2.250 1.100 2.845 1.475 ;
        RECT  1.750 0.325 2.250 1.475 ;
        RECT  1.100 0.325 1.750 0.690 ;
        RECT  1.100 1.100 1.750 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.780 0.740 0.890 ;
        RECT  0.250 0.700 0.350 1.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.165 3.200 0.165 ;
        RECT  2.960 -0.165 3.070 0.695 ;
        RECT  1.000 -0.165 2.960 0.165 ;
        RECT  0.870 -0.165 1.000 0.460 ;
        RECT  0.000 -0.165 0.870 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 1.635 3.200 1.965 ;
        RECT  2.960 1.050 3.070 1.965 ;
        RECT  0.990 1.635 2.960 1.965 ;
        RECT  0.880 1.260 0.990 1.965 ;
        RECT  0.000 1.635 0.880 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.325 2.850 0.690 ;
        RECT  2.350 1.100 2.845 1.475 ;
        RECT  1.100 0.325 1.650 0.690 ;
        RECT  1.100 1.100 1.650 1.475 ;
        RECT  2.495 0.800 2.925 0.940 ;
        RECT  0.990 0.800 1.590 0.940 ;
        RECT  0.850 0.570 0.990 1.150 ;
        RECT  0.740 0.570 0.850 0.690 ;
        RECT  0.740 1.030 0.850 1.150 ;
        RECT  0.610 0.295 0.740 0.690 ;
        RECT  0.610 1.030 0.740 1.470 ;
        RECT  0.050 0.435 0.610 0.545 ;
        RECT  0.050 1.245 0.610 1.355 ;
    END
END BUFFD8

MACRO BUFTD0
    CLASS CORE ;
    FOREIGN BUFTD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.310 1.950 1.490 ;
        RECT  1.820 0.310 1.850 0.490 ;
        RECT  1.820 1.255 1.850 1.490 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.105 ;
        RECT  1.150 1.005 1.250 1.105 ;
        RECT  1.050 1.005 1.150 1.490 ;
        RECT  0.550 1.400 1.050 1.490 ;
        RECT  0.450 1.055 0.550 1.490 ;
        RECT  0.350 1.055 0.450 1.145 ;
        RECT  0.250 0.775 0.350 1.145 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0565 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.895 ;
        RECT  0.955 0.725 1.050 0.895 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 -0.165 2.000 0.165 ;
        RECT  0.335 -0.165 0.445 0.455 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.875 1.760 0.985 ;
        RECT  1.640 0.320 1.730 0.765 ;
        RECT  0.800 0.320 1.640 0.420 ;
        RECT  1.440 0.510 1.530 1.455 ;
        RECT  1.295 0.510 1.440 0.600 ;
        RECT  1.275 1.345 1.440 1.455 ;
        RECT  0.800 1.055 0.940 1.225 ;
        RECT  0.700 0.320 0.800 1.225 ;
        RECT  0.555 0.320 0.700 0.420 ;
        RECT  0.500 0.565 0.600 0.935 ;
        RECT  0.180 0.565 0.500 0.665 ;
        RECT  0.160 0.275 0.180 0.665 ;
        RECT  0.160 1.255 0.180 1.490 ;
        RECT  0.070 0.275 0.160 1.490 ;
    END
END BUFTD0

MACRO BUFTD1
    CLASS CORE ;
    FOREIGN BUFTD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1200 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.310 1.950 1.490 ;
        RECT  1.820 0.310 1.850 0.490 ;
        RECT  1.820 1.110 1.850 1.490 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0832 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.105 ;
        RECT  1.150 1.005 1.250 1.105 ;
        RECT  1.050 1.005 1.150 1.490 ;
        RECT  0.550 1.400 1.050 1.490 ;
        RECT  0.450 1.055 0.550 1.490 ;
        RECT  0.350 1.055 0.450 1.145 ;
        RECT  0.250 0.775 0.350 1.145 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0839 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.895 ;
        RECT  0.955 0.725 1.050 0.895 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 -0.165 2.000 0.165 ;
        RECT  0.335 -0.165 0.445 0.455 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.895 1.760 1.005 ;
        RECT  1.640 0.320 1.730 0.785 ;
        RECT  0.800 0.320 1.640 0.420 ;
        RECT  1.440 0.510 1.530 1.455 ;
        RECT  1.295 0.510 1.440 0.600 ;
        RECT  1.275 1.345 1.440 1.455 ;
        RECT  0.800 1.055 0.940 1.225 ;
        RECT  0.700 0.320 0.800 1.225 ;
        RECT  0.555 0.320 0.700 0.420 ;
        RECT  0.500 0.565 0.600 0.935 ;
        RECT  0.180 0.565 0.500 0.665 ;
        RECT  0.160 0.275 0.180 0.665 ;
        RECT  0.160 1.255 0.180 1.490 ;
        RECT  0.070 0.275 0.160 1.490 ;
    END
END BUFTD1

MACRO BUFTD12
    CLASS CORE ;
    FOREIGN BUFTD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.9800 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.325 5.305 0.625 ;
        RECT  4.050 1.100 5.305 1.475 ;
        RECT  3.550 0.325 4.050 1.475 ;
        RECT  2.900 0.325 3.550 0.625 ;
        RECT  2.515 1.110 3.550 1.475 ;
        RECT  2.515 0.325 2.900 0.495 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.710 1.950 1.090 ;
        RECT  1.350 1.000 1.830 1.090 ;
        RECT  1.250 1.000 1.350 1.490 ;
        RECT  0.550 1.400 1.250 1.490 ;
        RECT  0.450 0.710 0.550 1.490 ;
        RECT  0.240 0.710 0.450 0.895 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1996 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.360 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.525 -0.165 5.600 0.165 ;
        RECT  5.415 -0.165 5.525 0.490 ;
        RECT  0.000 -0.165 5.415 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.525 1.635 5.600 1.965 ;
        RECT  5.415 1.110 5.525 1.965 ;
        RECT  0.000 1.635 5.415 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.150 0.325 5.305 0.625 ;
        RECT  4.150 1.100 5.305 1.475 ;
        RECT  2.900 0.325 3.450 0.625 ;
        RECT  2.515 1.110 3.450 1.475 ;
        RECT  2.515 0.325 2.900 0.495 ;
        RECT  2.415 0.650 2.710 0.770 ;
        RECT  2.185 0.880 2.710 1.000 ;
        RECT  2.275 0.305 2.415 0.770 ;
        RECT  1.140 0.305 2.275 0.420 ;
        RECT  2.055 0.510 2.185 1.385 ;
        RECT  1.775 0.510 2.055 0.620 ;
        RECT  1.505 1.230 2.055 1.385 ;
        RECT  1.050 0.305 1.140 1.250 ;
        RECT  0.525 0.305 1.050 0.420 ;
        RECT  0.765 1.150 1.050 1.250 ;
        RECT  0.850 0.510 0.950 0.920 ;
        RECT  0.175 0.510 0.850 0.600 ;
        RECT  0.150 0.310 0.175 0.600 ;
        RECT  0.150 1.065 0.175 1.490 ;
        RECT  0.060 0.310 0.150 1.490 ;
    END
END BUFTD12

MACRO BUFTD16
    CLASS CORE ;
    FOREIGN BUFTD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.3120 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.325 6.305 0.690 ;
        RECT  4.650 1.100 6.305 1.475 ;
        RECT  4.150 0.325 4.650 1.475 ;
        RECT  2.840 0.325 4.150 0.690 ;
        RECT  2.515 1.100 4.150 1.475 ;
        RECT  2.515 0.325 2.840 0.505 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.710 1.950 1.090 ;
        RECT  1.350 1.000 1.830 1.090 ;
        RECT  1.250 1.000 1.350 1.490 ;
        RECT  0.550 1.400 1.250 1.490 ;
        RECT  0.450 0.710 0.550 1.490 ;
        RECT  0.240 0.710 0.450 0.895 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1996 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.360 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.525 -0.165 6.600 0.165 ;
        RECT  6.415 -0.165 6.525 0.490 ;
        RECT  0.000 -0.165 6.415 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.525 1.635 6.600 1.965 ;
        RECT  6.415 1.110 6.525 1.965 ;
        RECT  0.000 1.635 6.415 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.750 0.325 6.305 0.690 ;
        RECT  4.750 1.100 6.305 1.475 ;
        RECT  2.840 0.325 4.050 0.690 ;
        RECT  2.515 1.100 4.050 1.475 ;
        RECT  2.515 0.325 2.840 0.505 ;
        RECT  2.425 0.615 2.710 0.750 ;
        RECT  2.195 0.870 2.710 1.000 ;
        RECT  2.285 0.280 2.425 0.750 ;
        RECT  1.140 0.280 2.285 0.420 ;
        RECT  2.055 0.510 2.195 1.385 ;
        RECT  1.765 0.510 2.055 0.620 ;
        RECT  1.505 1.215 2.055 1.385 ;
        RECT  1.050 0.280 1.140 1.250 ;
        RECT  0.525 0.280 1.050 0.420 ;
        RECT  0.765 1.150 1.050 1.250 ;
        RECT  0.850 0.510 0.950 0.920 ;
        RECT  0.175 0.510 0.850 0.600 ;
        RECT  0.150 0.310 0.175 0.600 ;
        RECT  0.150 1.065 0.175 1.490 ;
        RECT  0.060 0.310 0.150 1.490 ;
    END
END BUFTD16

MACRO BUFTD2
    CLASS CORE ;
    FOREIGN BUFTD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.825 0.310 1.950 1.490 ;
        RECT  1.770 0.310 1.825 0.555 ;
        RECT  1.760 1.115 1.825 1.490 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0803 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 0.710 1.300 1.155 ;
        RECT  1.100 1.055 1.200 1.155 ;
        RECT  1.000 1.055 1.100 1.490 ;
        RECT  0.550 1.400 1.000 1.490 ;
        RECT  0.450 1.055 0.550 1.490 ;
        RECT  0.340 1.055 0.450 1.145 ;
        RECT  0.230 0.775 0.340 1.145 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0769 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.510 0.965 0.920 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.200 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 0.895 1.710 1.005 ;
        RECT  1.590 0.275 1.680 0.785 ;
        RECT  0.750 0.275 1.590 0.375 ;
        RECT  1.390 0.510 1.480 1.455 ;
        RECT  1.240 0.510 1.390 0.600 ;
        RECT  1.215 1.345 1.390 1.455 ;
        RECT  0.750 1.100 0.890 1.275 ;
        RECT  0.660 0.275 0.750 1.275 ;
        RECT  0.525 0.275 0.660 0.420 ;
        RECT  0.460 0.565 0.570 0.860 ;
        RECT  0.180 0.565 0.460 0.665 ;
        RECT  0.140 0.330 0.180 0.665 ;
        RECT  0.140 1.255 0.180 1.490 ;
        RECT  0.050 0.330 0.140 1.490 ;
    END
END BUFTD2

MACRO BUFTD20
    CLASS CORE ;
    FOREIGN BUFTD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.6440 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.325 8.515 0.690 ;
        RECT  6.250 1.100 8.515 1.475 ;
        RECT  5.750 0.325 6.250 1.475 ;
        RECT  4.160 0.325 5.750 0.690 ;
        RECT  4.130 1.115 5.750 1.475 ;
        RECT  3.870 0.325 4.160 0.540 ;
        RECT  3.815 1.125 4.130 1.475 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1994 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.710 3.385 1.090 ;
        RECT  2.550 1.000 3.250 1.090 ;
        RECT  2.450 0.710 2.550 1.090 ;
        RECT  2.130 1.000 2.450 1.090 ;
        RECT  2.040 1.000 2.130 1.490 ;
        RECT  0.550 1.400 2.040 1.490 ;
        RECT  0.450 0.710 0.550 1.490 ;
        RECT  0.240 0.710 0.450 0.895 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.3048 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.760 1.090 ;
        RECT  0.950 1.000 1.650 1.090 ;
        RECT  0.850 0.710 0.950 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 8.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.635 8.800 1.965 ;
        RECT  3.500 1.450 3.690 1.965 ;
        RECT  0.000 1.635 3.500 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.350 0.325 8.515 0.690 ;
        RECT  6.350 1.100 8.515 1.475 ;
        RECT  4.130 1.115 5.650 1.475 ;
        RECT  3.870 0.325 4.160 0.540 ;
        RECT  3.815 1.125 4.130 1.475 ;
        RECT  3.780 0.640 4.020 0.775 ;
        RECT  3.585 0.870 4.020 1.015 ;
        RECT  3.675 0.280 3.780 0.775 ;
        RECT  1.950 0.280 3.675 0.420 ;
        RECT  3.475 0.510 3.585 1.340 ;
        RECT  2.330 0.510 3.475 0.620 ;
        RECT  2.355 1.200 3.475 1.340 ;
        RECT  2.220 1.200 2.355 1.470 ;
        RECT  1.850 0.280 1.950 1.300 ;
        RECT  0.525 0.280 1.850 0.420 ;
        RECT  0.735 1.200 1.850 1.300 ;
        RECT  1.250 0.510 1.350 0.885 ;
        RECT  0.175 0.510 1.250 0.600 ;
        RECT  0.150 0.310 0.175 0.600 ;
        RECT  0.150 1.065 0.175 1.490 ;
        RECT  0.060 0.310 0.150 1.490 ;
        RECT  4.160 0.325 5.650 0.690 ;
    END
END BUFTD20

MACRO BUFTD24
    CLASS CORE ;
    FOREIGN BUFTD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.9760 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.325 9.515 0.690 ;
        RECT  6.850 1.100 9.515 1.475 ;
        RECT  6.350 0.325 6.850 1.475 ;
        RECT  4.160 0.325 6.350 0.690 ;
        RECT  3.815 1.100 6.350 1.475 ;
        RECT  3.870 0.325 4.160 0.540 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1994 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.710 3.385 1.090 ;
        RECT  2.550 1.000 3.250 1.090 ;
        RECT  2.450 0.710 2.550 1.090 ;
        RECT  2.130 1.000 2.450 1.090 ;
        RECT  2.040 1.000 2.130 1.490 ;
        RECT  0.550 1.400 2.040 1.490 ;
        RECT  0.450 0.710 0.550 1.490 ;
        RECT  0.240 0.710 0.450 0.895 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.3048 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.760 1.090 ;
        RECT  0.950 1.000 1.650 1.090 ;
        RECT  0.850 0.710 0.950 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 9.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.635 9.800 1.965 ;
        RECT  3.500 1.430 3.690 1.965 ;
        RECT  0.000 1.635 3.500 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.950 0.325 9.515 0.690 ;
        RECT  4.160 0.325 6.250 0.690 ;
        RECT  3.815 1.100 6.250 1.475 ;
        RECT  3.870 0.325 4.160 0.540 ;
        RECT  3.780 0.640 4.020 0.780 ;
        RECT  3.580 0.870 4.020 1.000 ;
        RECT  3.670 0.280 3.780 0.780 ;
        RECT  1.950 0.280 3.670 0.420 ;
        RECT  3.475 0.510 3.580 1.340 ;
        RECT  2.330 0.510 3.475 0.620 ;
        RECT  2.330 1.200 3.475 1.340 ;
        RECT  2.220 1.200 2.330 1.470 ;
        RECT  1.850 0.280 1.950 1.300 ;
        RECT  0.525 0.280 1.850 0.420 ;
        RECT  0.735 1.200 1.850 1.300 ;
        RECT  1.250 0.510 1.350 0.885 ;
        RECT  0.175 0.510 1.250 0.600 ;
        RECT  0.150 0.330 0.175 0.600 ;
        RECT  0.150 1.065 0.175 1.490 ;
        RECT  0.060 0.330 0.150 1.490 ;
        RECT  6.950 1.100 9.515 1.475 ;
    END
END BUFTD24

MACRO BUFTD3
    CLASS CORE ;
    FOREIGN BUFTD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3120 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.310 2.485 0.490 ;
        RECT  2.250 1.110 2.485 1.490 ;
        RECT  1.950 0.310 2.250 1.490 ;
        RECT  1.820 0.310 1.950 0.490 ;
        RECT  1.820 1.110 1.950 1.490 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0832 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.105 ;
        RECT  1.150 1.005 1.250 1.105 ;
        RECT  1.050 1.005 1.150 1.490 ;
        RECT  0.550 1.400 1.050 1.490 ;
        RECT  0.450 1.055 0.550 1.490 ;
        RECT  0.350 1.055 0.450 1.145 ;
        RECT  0.250 0.775 0.350 1.145 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0839 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.895 ;
        RECT  0.955 0.725 1.050 0.895 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 -0.165 2.600 0.165 ;
        RECT  0.335 -0.165 0.445 0.455 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.310 2.485 0.490 ;
        RECT  2.350 1.110 2.485 1.490 ;
        RECT  1.820 0.310 1.850 0.490 ;
        RECT  1.820 1.110 1.850 1.490 ;
        RECT  1.730 0.645 1.830 0.755 ;
        RECT  1.530 0.895 1.760 1.005 ;
        RECT  1.640 0.320 1.730 0.755 ;
        RECT  0.800 0.320 1.640 0.420 ;
        RECT  1.440 0.510 1.530 1.455 ;
        RECT  1.295 0.510 1.440 0.600 ;
        RECT  1.275 1.345 1.440 1.455 ;
        RECT  0.800 1.055 0.940 1.225 ;
        RECT  0.700 0.320 0.800 1.225 ;
        RECT  0.555 0.320 0.700 0.420 ;
        RECT  0.500 0.565 0.600 0.935 ;
        RECT  0.180 0.565 0.500 0.665 ;
        RECT  0.160 0.275 0.180 0.665 ;
        RECT  0.160 1.255 0.180 1.490 ;
        RECT  0.070 0.275 0.160 1.490 ;
    END
END BUFTD3

MACRO BUFTD4
    CLASS CORE ;
    FOREIGN BUFTD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3160 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.310 2.485 0.490 ;
        RECT  2.250 1.110 2.485 1.490 ;
        RECT  1.950 0.310 2.250 1.490 ;
        RECT  1.820 0.310 1.950 0.490 ;
        RECT  1.820 1.110 1.950 1.490 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0832 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.105 ;
        RECT  1.150 1.005 1.250 1.105 ;
        RECT  1.050 1.005 1.150 1.490 ;
        RECT  0.550 1.400 1.050 1.490 ;
        RECT  0.450 1.055 0.550 1.490 ;
        RECT  0.350 1.055 0.450 1.145 ;
        RECT  0.250 0.775 0.350 1.145 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0839 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.895 ;
        RECT  0.910 0.725 1.050 0.895 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.705 -0.165 2.800 0.165 ;
        RECT  2.595 -0.165 2.705 0.550 ;
        RECT  0.445 -0.165 2.595 0.165 ;
        RECT  0.335 -0.165 0.445 0.455 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.705 1.635 2.800 1.965 ;
        RECT  2.595 1.110 2.705 1.965 ;
        RECT  0.000 1.635 2.595 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.310 2.485 0.490 ;
        RECT  2.350 1.110 2.485 1.490 ;
        RECT  1.820 0.310 1.850 0.490 ;
        RECT  1.820 1.110 1.850 1.490 ;
        RECT  1.730 0.645 1.830 0.755 ;
        RECT  1.530 0.895 1.760 1.005 ;
        RECT  1.640 0.320 1.730 0.755 ;
        RECT  0.800 0.320 1.640 0.420 ;
        RECT  1.440 0.510 1.530 1.455 ;
        RECT  1.295 0.510 1.440 0.600 ;
        RECT  1.275 1.345 1.440 1.455 ;
        RECT  0.800 1.055 0.940 1.225 ;
        RECT  0.700 0.320 0.800 1.225 ;
        RECT  0.555 0.320 0.700 0.420 ;
        RECT  0.500 0.565 0.600 0.935 ;
        RECT  0.180 0.565 0.500 0.665 ;
        RECT  0.160 0.275 0.180 0.665 ;
        RECT  0.160 1.255 0.180 1.490 ;
        RECT  0.070 0.275 0.160 1.490 ;
    END
END BUFTD4

MACRO BUFTD6
    CLASS CORE ;
    FOREIGN BUFTD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4820 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.310 3.705 0.490 ;
        RECT  3.250 1.110 3.705 1.490 ;
        RECT  2.950 0.310 3.250 1.490 ;
        RECT  2.515 0.310 2.950 0.490 ;
        RECT  2.515 1.110 2.950 1.490 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 1.950 1.090 ;
        RECT  1.350 1.000 1.850 1.090 ;
        RECT  1.250 1.000 1.350 1.490 ;
        RECT  0.550 1.400 1.250 1.490 ;
        RECT  0.450 0.710 0.550 1.490 ;
        RECT  0.240 0.710 0.450 0.895 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1996 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.360 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.925 -0.165 4.000 0.165 ;
        RECT  3.815 -0.165 3.925 0.560 ;
        RECT  0.000 -0.165 3.815 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.925 1.635 4.000 1.965 ;
        RECT  3.815 1.110 3.925 1.965 ;
        RECT  0.000 1.635 3.815 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.350 0.310 3.705 0.490 ;
        RECT  3.350 1.110 3.705 1.490 ;
        RECT  2.515 0.310 2.850 0.490 ;
        RECT  2.515 1.110 2.850 1.490 ;
        RECT  2.345 0.650 2.630 0.750 ;
        RECT  2.145 0.900 2.630 1.000 ;
        RECT  2.255 0.320 2.345 0.750 ;
        RECT  1.140 0.320 2.255 0.420 ;
        RECT  2.145 1.230 2.215 1.330 ;
        RECT  2.055 0.510 2.145 1.330 ;
        RECT  1.775 0.510 2.055 0.600 ;
        RECT  1.505 1.230 2.055 1.330 ;
        RECT  1.050 0.320 1.140 1.250 ;
        RECT  0.525 0.320 1.050 0.420 ;
        RECT  0.765 1.150 1.050 1.250 ;
        RECT  0.850 0.510 0.950 0.920 ;
        RECT  0.175 0.510 0.850 0.600 ;
        RECT  0.150 0.310 0.175 0.600 ;
        RECT  0.150 1.065 0.175 1.490 ;
        RECT  0.060 0.310 0.150 1.490 ;
    END
END BUFTD6

MACRO BUFTD8
    CLASS CORE ;
    FOREIGN BUFTD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.6480 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.325 4.305 0.690 ;
        RECT  3.650 1.100 4.305 1.475 ;
        RECT  3.150 0.325 3.650 1.475 ;
        RECT  2.890 0.325 3.150 0.690 ;
        RECT  2.555 1.130 3.150 1.475 ;
        RECT  2.555 0.325 2.890 0.540 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.710 1.950 1.090 ;
        RECT  1.350 1.000 1.830 1.090 ;
        RECT  1.250 1.000 1.350 1.490 ;
        RECT  0.550 1.400 1.250 1.490 ;
        RECT  0.450 0.710 0.550 1.490 ;
        RECT  0.240 0.710 0.450 0.895 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1993 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.360 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 -0.165 4.600 0.165 ;
        RECT  4.415 -0.165 4.525 0.490 ;
        RECT  0.000 -0.165 4.415 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.635 4.600 1.965 ;
        RECT  4.415 1.110 4.525 1.965 ;
        RECT  2.435 1.635 4.415 1.965 ;
        RECT  2.325 1.130 2.435 1.965 ;
        RECT  0.000 1.635 2.325 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 0.325 4.305 0.690 ;
        RECT  3.750 1.100 4.305 1.475 ;
        RECT  2.890 0.325 3.050 0.690 ;
        RECT  2.555 1.130 3.050 1.475 ;
        RECT  2.555 0.325 2.890 0.540 ;
        RECT  2.465 0.650 2.750 0.780 ;
        RECT  2.215 0.870 2.750 1.020 ;
        RECT  2.325 0.280 2.465 0.780 ;
        RECT  1.140 0.280 2.325 0.420 ;
        RECT  2.075 0.510 2.215 1.370 ;
        RECT  1.765 0.510 2.075 0.620 ;
        RECT  1.505 1.230 2.075 1.370 ;
        RECT  1.050 0.280 1.140 1.250 ;
        RECT  0.525 0.280 1.050 0.420 ;
        RECT  0.765 1.125 1.050 1.250 ;
        RECT  0.850 0.510 0.950 0.920 ;
        RECT  0.175 0.510 0.850 0.600 ;
        RECT  0.150 0.310 0.175 0.600 ;
        RECT  0.150 1.065 0.175 1.490 ;
        RECT  0.060 0.310 0.150 1.490 ;
    END
END BUFTD8

MACRO CKAN2D0
    CLASS CORE ;
    FOREIGN CKAN2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.460 1.150 1.090 ;
        RECT  0.900 0.460 1.050 0.570 ;
        RECT  1.040 0.980 1.050 1.090 ;
        RECT  0.930 0.980 1.040 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0214 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.575 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0207 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.210 0.710 0.250 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.805 -0.165 1.200 0.165 ;
        RECT  0.635 -0.165 0.805 0.370 ;
        RECT  0.000 -0.165 0.635 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.635 1.200 1.965 ;
        RECT  0.615 1.390 0.820 1.965 ;
        RECT  0.230 1.635 0.615 1.965 ;
        RECT  0.120 1.205 0.230 1.965 ;
        RECT  0.000 1.635 0.120 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.785 0.780 0.935 0.890 ;
        RECT  0.685 0.460 0.785 1.300 ;
        RECT  0.070 0.460 0.685 0.570 ;
        RECT  0.330 1.210 0.685 1.300 ;
    END
END CKAN2D0

MACRO CKAN2D1
    CLASS CORE ;
    FOREIGN CKAN2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.465 1.150 1.090 ;
        RECT  0.900 0.465 1.050 0.575 ;
        RECT  1.040 0.980 1.050 1.090 ;
        RECT  0.930 0.980 1.040 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0244 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.575 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.210 0.710 0.250 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.805 -0.165 1.200 0.165 ;
        RECT  0.635 -0.165 0.805 0.370 ;
        RECT  0.000 -0.165 0.635 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.635 1.200 1.965 ;
        RECT  0.615 1.390 0.820 1.965 ;
        RECT  0.230 1.635 0.615 1.965 ;
        RECT  0.120 1.205 0.230 1.965 ;
        RECT  0.000 1.635 0.120 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.785 0.780 0.935 0.890 ;
        RECT  0.685 0.460 0.785 1.300 ;
        RECT  0.070 0.460 0.685 0.570 ;
        RECT  0.330 1.210 0.685 1.300 ;
    END
END CKAN2D1

MACRO CKAN2D2
    CLASS CORE ;
    FOREIGN CKAN2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1780 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.275 1.150 1.495 ;
        RECT  0.940 0.275 1.050 0.675 ;
        RECT  0.900 1.390 1.050 1.495 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0438 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.570 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.350 1.100 ;
        RECT  0.200 0.700 0.250 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.795 -0.165 1.400 0.165 ;
        RECT  0.625 -0.165 0.795 0.350 ;
        RECT  0.000 -0.165 0.625 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.635 1.400 1.965 ;
        RECT  0.630 1.410 0.790 1.965 ;
        RECT  0.220 1.635 0.630 1.965 ;
        RECT  0.110 1.210 0.220 1.965 ;
        RECT  0.000 1.635 0.110 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.460 0.830 1.300 ;
        RECT  0.065 0.460 0.720 0.570 ;
        RECT  0.485 1.210 0.720 1.300 ;
        RECT  0.375 1.210 0.485 1.420 ;
    END
END CKAN2D2

MACRO CKAN2D4
    CLASS CORE ;
    FOREIGN CKAN2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.390 1.515 1.495 ;
        RECT  1.150 0.310 1.450 1.495 ;
        RECT  0.940 0.310 1.150 0.690 ;
        RECT  0.795 1.390 1.150 1.495 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0438 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.570 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.350 1.100 ;
        RECT  0.195 0.700 0.250 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.795 -0.165 1.800 0.165 ;
        RECT  0.625 -0.165 0.795 0.350 ;
        RECT  0.000 -0.165 0.625 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.620 1.030 1.725 1.965 ;
        RECT  0.185 1.635 1.620 1.965 ;
        RECT  0.075 1.210 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 0.310 1.050 0.690 ;
        RECT  0.795 1.390 1.050 1.495 ;
        RECT  0.720 0.460 0.830 1.300 ;
        RECT  0.065 0.460 0.720 0.570 ;
        RECT  0.450 1.210 0.720 1.300 ;
        RECT  0.335 1.210 0.450 1.420 ;
    END
END CKAN2D4

MACRO CKAN2D8
    CLASS CORE ;
    FOREIGN CKAN2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.5760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.115 3.105 1.475 ;
        RECT  2.250 0.325 3.080 0.690 ;
        RECT  1.750 0.325 2.250 1.475 ;
        RECT  1.395 0.325 1.750 0.690 ;
        RECT  1.395 1.105 1.750 1.475 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0708 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.710 1.065 0.940 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.350 1.000 0.850 1.090 ;
        RECT  0.245 0.710 0.350 1.090 ;
        RECT  0.175 0.710 0.245 0.945 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0702 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.335 -0.165 3.400 0.165 ;
        RECT  3.205 -0.165 3.335 0.495 ;
        RECT  0.215 -0.165 3.205 0.165 ;
        RECT  0.085 -0.165 0.215 0.495 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.325 1.635 3.400 1.965 ;
        RECT  3.215 1.050 3.325 1.965 ;
        RECT  0.970 1.635 3.215 1.965 ;
        RECT  0.970 1.400 1.285 1.510 ;
        RECT  0.830 1.400 0.970 1.965 ;
        RECT  0.560 1.400 0.830 1.510 ;
        RECT  0.205 1.635 0.830 1.965 ;
        RECT  0.095 1.215 0.205 1.965 ;
        RECT  0.000 1.635 0.095 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 1.115 3.105 1.475 ;
        RECT  2.350 0.325 3.080 0.690 ;
        RECT  1.395 0.325 1.650 0.690 ;
        RECT  1.395 1.105 1.650 1.475 ;
        RECT  2.410 0.800 3.170 0.940 ;
        RECT  1.305 0.800 1.590 0.940 ;
        RECT  1.165 0.335 1.305 1.310 ;
        RECT  0.565 0.335 1.165 0.475 ;
        RECT  0.315 1.180 1.165 1.310 ;
    END
END CKAN2D8

MACRO CKBD0
    CLASS CORE ;
    FOREIGN CKBD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.275 0.750 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0246 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 -0.165 0.800 0.165 ;
        RECT  0.295 -0.165 0.495 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 1.635 0.800 1.965 ;
        RECT  0.335 1.260 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.445 0.510 0.535 1.150 ;
        RECT  0.185 0.510 0.445 0.600 ;
        RECT  0.185 1.040 0.445 1.150 ;
        RECT  0.075 0.275 0.185 0.600 ;
        RECT  0.075 1.040 0.185 1.490 ;
    END
END CKBD0

MACRO CKBD1
    CLASS CORE ;
    FOREIGN CKBD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1330 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.310 0.750 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 -0.165 0.800 0.165 ;
        RECT  0.305 -0.165 0.495 0.400 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 1.635 0.800 1.965 ;
        RECT  0.345 1.260 0.455 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.445 0.510 0.535 1.150 ;
        RECT  0.185 0.510 0.445 0.600 ;
        RECT  0.185 1.040 0.445 1.150 ;
        RECT  0.075 0.310 0.185 0.600 ;
        RECT  0.075 1.040 0.185 1.470 ;
    END
END CKBD1

MACRO CKBD12
    CLASS CORE ;
    FOREIGN CKBD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.0050 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.100 4.100 1.475 ;
        RECT  2.850 0.325 3.645 0.690 ;
        RECT  2.350 0.325 2.850 1.475 ;
        RECT  1.375 0.325 2.350 0.690 ;
        RECT  1.310 1.100 2.350 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1966 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.775 0.710 0.925 ;
        RECT  0.050 0.275 0.210 0.925 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.875 -0.165 4.400 0.165 ;
        RECT  3.745 -0.165 3.875 0.495 ;
        RECT  1.260 -0.165 3.745 0.165 ;
        RECT  1.130 -0.165 1.260 0.690 ;
        RECT  0.000 -0.165 1.130 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.320 1.635 4.400 1.965 ;
        RECT  4.210 1.050 4.320 1.965 ;
        RECT  1.210 1.635 4.210 1.965 ;
        RECT  1.080 1.030 1.210 1.965 ;
        RECT  0.000 1.635 1.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 1.100 4.100 1.475 ;
        RECT  2.950 0.325 3.645 0.690 ;
        RECT  1.375 0.325 2.250 0.690 ;
        RECT  1.310 1.100 2.250 1.475 ;
        RECT  3.010 0.800 4.155 0.940 ;
        RECT  0.980 0.800 2.140 0.940 ;
        RECT  0.840 0.275 0.980 1.500 ;
        RECT  0.480 0.545 0.840 0.685 ;
        RECT  0.820 1.040 0.840 1.500 ;
        RECT  0.450 1.040 0.820 1.180 ;
        RECT  0.350 0.275 0.480 0.685 ;
        RECT  0.320 1.040 0.450 1.500 ;
    END
END CKBD12

MACRO CKBD16
    CLASS CORE ;
    FOREIGN CKBD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.3490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.110 5.305 1.475 ;
        RECT  3.450 0.325 4.970 0.690 ;
        RECT  2.950 0.325 3.450 1.475 ;
        RECT  1.660 0.325 2.950 0.690 ;
        RECT  1.565 1.110 2.950 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2516 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.220 0.790 0.950 0.910 ;
        RECT  0.050 0.275 0.220 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.550 -0.165 5.600 0.165 ;
        RECT  1.415 -0.165 1.550 0.690 ;
        RECT  0.515 -0.165 1.415 0.165 ;
        RECT  0.385 -0.165 0.515 0.680 ;
        RECT  0.000 -0.165 0.385 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.525 1.635 5.600 1.965 ;
        RECT  5.415 1.040 5.525 1.965 ;
        RECT  0.000 1.635 5.415 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.550 1.110 5.305 1.475 ;
        RECT  3.550 0.325 4.970 0.690 ;
        RECT  1.660 0.325 2.850 0.690 ;
        RECT  1.565 1.110 2.850 1.475 ;
        RECT  3.620 0.800 5.205 0.940 ;
        RECT  1.295 0.800 2.790 0.940 ;
        RECT  1.125 0.285 1.295 1.500 ;
        RECT  1.090 0.510 1.125 1.500 ;
        RECT  0.775 0.510 1.090 0.680 ;
        RECT  0.705 1.040 1.090 1.210 ;
        RECT  0.645 0.275 0.775 0.680 ;
        RECT  0.575 1.040 0.705 1.500 ;
        RECT  0.190 1.040 0.575 1.210 ;
        RECT  0.070 1.040 0.190 1.500 ;
    END
END CKBD16

MACRO CKBD2
    CLASS CORE ;
    FOREIGN CKBD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1660 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 0.560 1.150 1.150 ;
        RECT  0.865 0.560 1.025 0.670 ;
        RECT  0.865 1.020 1.025 1.150 ;
        RECT  0.755 0.310 0.865 0.670 ;
        RECT  0.755 1.020 0.865 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.710 0.365 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.125 -0.165 1.200 0.165 ;
        RECT  1.015 -0.165 1.125 0.450 ;
        RECT  0.640 -0.165 1.015 0.165 ;
        RECT  0.465 -0.165 0.640 0.400 ;
        RECT  0.000 -0.165 0.465 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.125 1.635 1.200 1.965 ;
        RECT  1.015 1.260 1.125 1.965 ;
        RECT  0.610 1.635 1.015 1.965 ;
        RECT  0.485 1.260 0.610 1.965 ;
        RECT  0.000 1.635 0.485 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 0.780 0.850 0.890 ;
        RECT  0.600 0.490 0.605 0.890 ;
        RECT  0.495 0.490 0.600 1.120 ;
        RECT  0.345 0.490 0.495 0.600 ;
        RECT  0.345 1.030 0.495 1.120 ;
        RECT  0.235 0.310 0.345 0.600 ;
        RECT  0.235 1.030 0.345 1.470 ;
    END
END CKBD2

MACRO CKBD20
    CLASS CORE ;
    FOREIGN CKBD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.6600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 1.100 6.505 1.475 ;
        RECT  4.050 0.325 5.730 0.690 ;
        RECT  3.550 0.325 4.050 1.475 ;
        RECT  1.910 0.325 3.550 0.690 ;
        RECT  1.795 1.100 3.550 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3003 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 0.805 1.200 0.920 ;
        RECT  0.050 0.275 0.190 0.920 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.960 -0.165 6.800 0.165 ;
        RECT  5.850 -0.165 5.960 0.495 ;
        RECT  1.785 -0.165 5.850 0.165 ;
        RECT  1.675 -0.165 1.785 0.695 ;
        RECT  0.000 -0.165 1.675 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 1.635 6.800 1.965 ;
        RECT  6.615 1.040 6.725 1.965 ;
        RECT  0.185 1.635 6.615 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.150 1.100 6.505 1.475 ;
        RECT  4.150 0.325 5.730 0.690 ;
        RECT  1.910 0.325 3.450 0.690 ;
        RECT  1.795 1.100 3.450 1.475 ;
        RECT  4.210 0.800 6.480 0.940 ;
        RECT  1.550 0.800 3.365 0.940 ;
        RECT  1.350 0.280 1.550 1.505 ;
        RECT  1.335 0.475 1.350 1.505 ;
        RECT  0.985 0.475 1.335 0.675 ;
        RECT  0.955 1.045 1.335 1.245 ;
        RECT  0.875 0.280 0.985 0.675 ;
        RECT  0.825 1.045 0.955 1.505 ;
        RECT  0.465 0.475 0.875 0.675 ;
        RECT  0.455 1.045 0.825 1.245 ;
        RECT  0.355 0.280 0.465 0.675 ;
        RECT  0.325 1.045 0.455 1.505 ;
    END
END CKBD20

MACRO CKBD24
    CLASS CORE ;
    FOREIGN CKBD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 2.0540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 1.100 7.735 1.475 ;
        RECT  4.850 0.325 7.480 0.670 ;
        RECT  4.350 0.325 4.850 1.475 ;
        RECT  2.090 0.325 4.350 0.670 ;
        RECT  2.045 1.100 4.350 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3487 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 0.805 1.260 0.920 ;
        RECT  0.050 0.275 0.190 0.920 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.975 -0.165 7.800 0.165 ;
        RECT  1.845 -0.165 1.975 0.665 ;
        RECT  0.000 -0.165 1.845 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 7.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.950 1.100 7.735 1.475 ;
        RECT  4.950 0.325 7.480 0.670 ;
        RECT  2.090 0.325 4.250 0.670 ;
        RECT  2.045 1.100 4.250 1.475 ;
        RECT  5.190 0.780 7.380 0.920 ;
        RECT  1.735 0.780 4.190 0.905 ;
        RECT  1.505 0.365 1.735 1.500 ;
        RECT  0.550 0.365 1.505 0.595 ;
        RECT  1.185 1.270 1.505 1.500 ;
        RECT  1.075 1.040 1.185 1.500 ;
        RECT  0.685 1.270 1.075 1.500 ;
        RECT  0.575 1.040 0.685 1.500 ;
        RECT  0.185 1.270 0.575 1.500 ;
        RECT  0.075 1.040 0.185 1.500 ;
    END
END CKBD24

MACRO CKBD3
    CLASS CORE ;
    FOREIGN CKBD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2990 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.340 1.350 0.590 ;
        RECT  1.250 1.060 1.350 1.490 ;
        RECT  1.200 0.340 1.250 1.490 ;
        RECT  0.950 0.340 1.200 1.250 ;
        RECT  0.695 0.340 0.950 0.590 ;
        RECT  0.815 1.060 0.950 1.250 ;
        RECT  0.695 1.060 0.815 1.470 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.710 0.355 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.165 1.400 0.165 ;
        RECT  0.405 -0.165 0.580 0.400 ;
        RECT  0.000 -0.165 0.405 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.565 1.635 1.400 1.965 ;
        RECT  0.425 1.260 0.565 1.965 ;
        RECT  0.000 1.635 0.425 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.695 0.340 0.850 0.590 ;
        RECT  0.815 1.060 0.850 1.250 ;
        RECT  0.695 1.060 0.815 1.470 ;
        RECT  0.565 0.780 0.790 0.890 ;
        RECT  0.545 0.490 0.565 0.890 ;
        RECT  0.445 0.490 0.545 1.120 ;
        RECT  0.285 0.490 0.445 0.600 ;
        RECT  0.285 1.030 0.445 1.120 ;
        RECT  0.175 0.310 0.285 0.600 ;
        RECT  0.175 1.030 0.285 1.470 ;
    END
END CKBD3

MACRO CKBD4
    CLASS CORE ;
    FOREIGN CKBD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.310 1.505 0.690 ;
        RECT  1.450 1.110 1.505 1.490 ;
        RECT  1.150 0.310 1.450 1.490 ;
        RECT  0.805 0.310 1.150 0.690 ;
        RECT  0.805 1.110 1.150 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1003 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.355 0.920 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.520 ;
        RECT  0.185 -0.165 1.615 0.165 ;
        RECT  0.075 -0.165 0.185 0.520 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.040 1.725 1.965 ;
        RECT  0.185 1.635 1.615 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.805 0.310 1.050 0.690 ;
        RECT  0.805 1.110 1.050 1.490 ;
        RECT  0.695 0.780 0.930 0.890 ;
        RECT  0.585 0.360 0.695 1.140 ;
        RECT  0.295 0.360 0.585 0.470 ;
        RECT  0.445 1.040 0.585 1.140 ;
        RECT  0.335 1.040 0.445 1.490 ;
    END
END CKBD4

MACRO CKBD6
    CLASS CORE ;
    FOREIGN CKBD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.5200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.310 2.305 0.690 ;
        RECT  1.650 1.110 2.045 1.490 ;
        RECT  1.350 0.310 1.650 1.490 ;
        RECT  1.080 0.310 1.350 0.690 ;
        RECT  0.815 1.110 1.350 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0948 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.510 0.355 0.920 ;
        RECT  0.185 0.510 0.245 0.705 ;
        RECT  0.050 0.275 0.185 0.705 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.960 -0.165 2.400 0.165 ;
        RECT  0.830 -0.165 0.960 0.510 ;
        RECT  0.000 -0.165 0.830 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.265 1.635 2.400 1.965 ;
        RECT  2.155 1.040 2.265 1.965 ;
        RECT  0.705 1.635 2.155 1.965 ;
        RECT  0.595 1.260 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.750 0.310 2.305 0.690 ;
        RECT  1.750 1.110 2.045 1.490 ;
        RECT  1.080 0.310 1.250 0.690 ;
        RECT  0.815 1.110 1.250 1.490 ;
        RECT  0.675 0.800 1.220 0.910 ;
        RECT  0.565 0.310 0.675 1.140 ;
        RECT  0.445 1.040 0.565 1.140 ;
        RECT  0.335 1.040 0.445 1.500 ;
    END
END CKBD6

MACRO CKBD8
    CLASS CORE ;
    FOREIGN CKBD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.6960 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.325 2.925 0.690 ;
        RECT  2.250 1.100 2.825 1.475 ;
        RECT  1.750 0.325 2.250 1.475 ;
        RECT  1.175 0.325 1.750 0.690 ;
        RECT  1.075 1.100 1.750 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1412 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.510 0.355 0.920 ;
        RECT  0.245 0.275 0.255 0.920 ;
        RECT  0.145 0.275 0.245 0.705 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.165 3.200 0.165 ;
        RECT  0.940 -0.165 1.050 0.695 ;
        RECT  0.000 -0.165 0.940 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.045 1.635 3.200 1.965 ;
        RECT  2.935 1.040 3.045 1.965 ;
        RECT  0.965 1.635 2.935 1.965 ;
        RECT  0.855 1.070 0.965 1.965 ;
        RECT  0.445 1.635 0.855 1.965 ;
        RECT  0.335 1.290 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.325 2.925 0.690 ;
        RECT  2.350 1.100 2.825 1.475 ;
        RECT  1.175 0.325 1.650 0.690 ;
        RECT  1.075 1.100 1.650 1.475 ;
        RECT  2.385 0.800 2.815 0.940 ;
        RECT  0.770 0.800 1.580 0.940 ;
        RECT  0.735 0.275 0.770 0.940 ;
        RECT  0.595 0.275 0.735 1.500 ;
        RECT  0.185 1.040 0.595 1.180 ;
        RECT  0.075 1.040 0.185 1.500 ;
    END
END CKBD8

MACRO CKLHQD1
    CLASS CORE ;
    FOREIGN CKLHQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.825 0.275 3.950 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0830 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.710 2.365 1.090 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.455 -0.165 4.000 0.165 ;
        RECT  1.285 -0.165 1.455 0.450 ;
        RECT  0.000 -0.165 1.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.635 4.000 1.965 ;
        RECT  1.280 1.445 1.490 1.965 ;
        RECT  0.185 1.635 1.280 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.595 0.740 3.695 1.490 ;
        RECT  2.710 1.400 3.595 1.490 ;
        RECT  3.385 0.465 3.475 1.155 ;
        RECT  3.340 0.465 3.385 0.655 ;
        RECT  3.045 1.055 3.385 1.155 ;
        RECT  3.245 0.760 3.295 0.940 ;
        RECT  3.145 0.275 3.245 0.940 ;
        RECT  1.755 0.275 3.145 0.365 ;
        RECT  2.945 0.740 3.045 1.155 ;
        RECT  2.710 0.505 2.985 0.615 ;
        RECT  2.600 0.505 2.710 1.490 ;
        RECT  2.115 0.505 2.510 0.615 ;
        RECT  2.115 1.310 2.475 1.420 ;
        RECT  2.025 0.505 2.115 1.420 ;
        RECT  1.845 0.475 1.935 1.515 ;
        RECT  1.825 1.265 1.845 1.515 ;
        RECT  1.150 1.265 1.825 1.355 ;
        RECT  1.665 0.275 1.755 1.155 ;
        RECT  1.545 0.275 1.665 0.465 ;
        RECT  1.295 1.055 1.665 1.155 ;
        RECT  1.450 0.560 1.550 0.940 ;
        RECT  1.070 0.560 1.450 0.660 ;
        RECT  1.195 0.750 1.295 1.155 ;
        RECT  1.050 1.265 1.150 1.495 ;
        RECT  0.970 0.315 1.070 1.155 ;
        RECT  0.740 1.385 1.050 1.495 ;
        RECT  0.805 0.315 0.970 0.425 ;
        RECT  0.940 1.055 0.970 1.155 ;
        RECT  0.830 1.055 0.940 1.295 ;
        RECT  0.740 0.555 0.880 0.665 ;
        RECT  0.640 0.555 0.740 1.495 ;
        RECT  0.185 0.315 0.715 0.425 ;
        RECT  0.075 0.315 0.185 0.565 ;
    END
END CKLHQD1

MACRO CKLHQD12
    CLASS CORE ;
    FOREIGN CKLHQD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.0920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.325 7.315 0.695 ;
        RECT  6.250 1.100 7.315 1.475 ;
        RECT  5.750 0.325 6.250 1.475 ;
        RECT  4.665 0.325 5.750 0.695 ;
        RECT  4.665 1.100 5.750 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.1768 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.190 0.710 4.320 1.295 ;
        RECT  3.355 1.205 4.190 1.295 ;
        RECT  3.245 0.710 3.355 1.295 ;
        RECT  2.355 1.205 3.245 1.295 ;
        RECT  2.245 0.710 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 7.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.945 1.635 7.600 1.965 ;
        RECT  2.755 1.390 2.945 1.965 ;
        RECT  1.475 1.635 2.755 1.965 ;
        RECT  1.265 1.445 1.475 1.965 ;
        RECT  0.185 1.635 1.265 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.350 0.325 7.315 0.695 ;
        RECT  6.350 1.100 7.315 1.475 ;
        RECT  4.665 0.325 5.650 0.695 ;
        RECT  4.665 1.100 5.650 1.475 ;
        RECT  6.430 0.805 7.300 0.945 ;
        RECT  4.575 0.805 5.575 0.945 ;
        RECT  4.435 0.300 4.575 1.525 ;
        RECT  3.025 0.300 4.435 0.440 ;
        RECT  3.215 1.385 4.435 1.525 ;
        RECT  3.750 0.530 3.850 0.895 ;
        RECT  3.040 0.530 3.750 0.620 ;
        RECT  2.950 0.530 3.040 1.115 ;
        RECT  2.670 1.025 2.950 1.115 ;
        RECT  2.570 0.475 2.670 1.115 ;
        RECT  1.700 0.275 2.570 0.365 ;
        RECT  2.500 1.025 2.570 1.115 ;
        RECT  2.120 1.390 2.470 1.490 ;
        RECT  2.120 0.505 2.460 0.615 ;
        RECT  2.030 0.505 2.120 1.490 ;
        RECT  1.970 0.835 2.030 1.025 ;
        RECT  1.880 0.505 1.940 0.715 ;
        RECT  1.880 1.265 1.920 1.515 ;
        RECT  1.820 0.505 1.880 1.515 ;
        RECT  1.790 0.505 1.820 1.355 ;
        RECT  1.150 1.265 1.790 1.355 ;
        RECT  1.610 0.275 1.700 1.155 ;
        RECT  1.525 0.275 1.610 0.450 ;
        RECT  1.295 1.055 1.610 1.155 ;
        RECT  1.400 0.545 1.500 0.785 ;
        RECT  1.070 0.545 1.400 0.635 ;
        RECT  1.195 0.885 1.295 1.155 ;
        RECT  1.050 1.265 1.150 1.495 ;
        RECT  0.970 0.315 1.070 1.155 ;
        RECT  0.740 1.385 1.050 1.495 ;
        RECT  0.805 0.315 0.970 0.425 ;
        RECT  0.940 1.055 0.970 1.155 ;
        RECT  0.830 1.055 0.940 1.295 ;
        RECT  0.740 0.555 0.880 0.665 ;
        RECT  0.640 0.555 0.740 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD12

MACRO CKLHQD16
    CLASS CORE ;
    FOREIGN CKLHQD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.4560 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.325 8.905 0.695 ;
        RECT  7.250 1.100 8.905 1.475 ;
        RECT  6.750 0.325 7.250 1.475 ;
        RECT  5.265 0.325 6.750 0.695 ;
        RECT  5.265 1.100 6.750 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.2489 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.710 4.555 1.295 ;
        RECT  3.555 1.205 4.445 1.295 ;
        RECT  3.445 0.710 3.555 1.295 ;
        RECT  2.355 1.205 3.445 1.295 ;
        RECT  2.245 0.710 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.125 -0.165 9.200 0.165 ;
        RECT  9.015 -0.165 9.125 0.690 ;
        RECT  0.000 -0.165 9.015 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.125 1.635 9.200 1.965 ;
        RECT  9.015 1.110 9.125 1.965 ;
        RECT  3.175 1.635 9.015 1.965 ;
        RECT  2.985 1.390 3.175 1.965 ;
        RECT  1.435 1.635 2.985 1.965 ;
        RECT  1.245 1.445 1.435 1.965 ;
        RECT  0.185 1.635 1.245 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.350 0.325 8.905 0.695 ;
        RECT  7.350 1.100 8.905 1.475 ;
        RECT  5.265 0.325 6.650 0.695 ;
        RECT  5.265 1.100 6.650 1.475 ;
        RECT  7.410 0.805 8.950 0.945 ;
        RECT  5.175 0.805 6.590 0.945 ;
        RECT  5.035 0.305 5.175 1.525 ;
        RECT  3.215 0.305 5.035 0.440 ;
        RECT  3.455 1.390 5.035 1.525 ;
        RECT  4.830 0.530 4.945 0.915 ;
        RECT  4.065 0.530 4.830 0.620 ;
        RECT  3.935 0.530 4.065 0.895 ;
        RECT  3.260 0.530 3.935 0.620 ;
        RECT  3.140 0.530 3.260 1.115 ;
        RECT  2.860 1.015 3.140 1.115 ;
        RECT  2.760 0.475 2.860 1.115 ;
        RECT  2.720 1.015 2.760 1.115 ;
        RECT  2.550 0.275 2.650 0.895 ;
        RECT  1.670 0.275 2.550 0.365 ;
        RECT  2.090 1.390 2.440 1.490 ;
        RECT  2.090 0.505 2.430 0.615 ;
        RECT  2.000 0.505 2.090 1.490 ;
        RECT  1.940 0.825 2.000 1.015 ;
        RECT  1.850 0.505 1.890 0.705 ;
        RECT  1.850 1.265 1.890 1.515 ;
        RECT  1.790 0.505 1.850 1.515 ;
        RECT  1.760 0.505 1.790 1.355 ;
        RECT  1.135 1.265 1.760 1.355 ;
        RECT  1.580 0.275 1.670 1.155 ;
        RECT  1.485 0.275 1.580 0.450 ;
        RECT  1.270 1.055 1.580 1.155 ;
        RECT  1.370 0.545 1.470 0.785 ;
        RECT  1.070 0.545 1.370 0.635 ;
        RECT  1.170 0.905 1.270 1.155 ;
        RECT  1.040 1.265 1.135 1.495 ;
        RECT  0.970 0.310 1.070 1.155 ;
        RECT  0.730 1.385 1.040 1.495 ;
        RECT  0.805 0.310 0.970 0.420 ;
        RECT  0.930 1.055 0.970 1.155 ;
        RECT  0.820 1.055 0.930 1.295 ;
        RECT  0.730 0.535 0.880 0.645 ;
        RECT  0.640 0.535 0.730 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD16

MACRO CKLHQD2
    CLASS CORE ;
    FOREIGN CKLHQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.865 0.545 3.950 1.205 ;
        RECT  3.850 0.275 3.865 1.490 ;
        RECT  3.755 0.275 3.850 0.675 ;
        RECT  3.755 1.055 3.850 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0830 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.710 2.355 1.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 -0.165 4.200 0.165 ;
        RECT  4.010 -0.165 4.130 0.455 ;
        RECT  0.000 -0.165 4.010 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 1.635 4.200 1.965 ;
        RECT  4.010 1.325 4.130 1.965 ;
        RECT  1.475 1.635 4.010 1.965 ;
        RECT  1.265 1.445 1.475 1.965 ;
        RECT  0.185 1.635 1.265 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.540 0.740 3.640 1.375 ;
        RECT  2.645 1.285 3.540 1.375 ;
        RECT  3.330 0.465 3.420 1.165 ;
        RECT  3.285 0.465 3.330 0.655 ;
        RECT  2.990 1.065 3.330 1.165 ;
        RECT  3.190 0.760 3.240 0.950 ;
        RECT  3.090 0.275 3.190 0.950 ;
        RECT  1.700 0.275 3.090 0.365 ;
        RECT  2.890 0.740 2.990 1.165 ;
        RECT  2.645 0.505 2.940 0.615 ;
        RECT  2.545 0.505 2.645 1.375 ;
        RECT  2.120 0.505 2.455 0.615 ;
        RECT  2.325 1.265 2.425 1.515 ;
        RECT  2.120 1.265 2.325 1.355 ;
        RECT  2.030 0.505 2.120 1.355 ;
        RECT  1.970 0.835 2.030 1.025 ;
        RECT  1.880 0.505 1.920 0.705 ;
        RECT  1.880 1.265 1.920 1.515 ;
        RECT  1.820 0.505 1.880 1.515 ;
        RECT  1.790 0.505 1.820 1.355 ;
        RECT  1.150 1.265 1.790 1.355 ;
        RECT  1.610 0.275 1.700 1.155 ;
        RECT  1.525 0.275 1.610 0.450 ;
        RECT  1.295 1.055 1.610 1.155 ;
        RECT  1.400 0.545 1.500 0.785 ;
        RECT  1.070 0.545 1.400 0.635 ;
        RECT  1.195 0.885 1.295 1.155 ;
        RECT  1.050 1.265 1.150 1.495 ;
        RECT  0.970 0.315 1.070 1.155 ;
        RECT  0.740 1.385 1.050 1.495 ;
        RECT  0.805 0.315 0.970 0.425 ;
        RECT  0.940 1.055 0.970 1.155 ;
        RECT  0.830 1.055 0.940 1.295 ;
        RECT  0.740 0.555 0.880 0.665 ;
        RECT  0.640 0.555 0.740 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD2

MACRO CKLHQD20
    CLASS CORE ;
    FOREIGN CKLHQD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.8200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.325 9.905 0.690 ;
        RECT  7.650 1.100 9.905 1.475 ;
        RECT  7.150 0.325 7.650 1.475 ;
        RECT  5.265 0.325 7.150 0.695 ;
        RECT  5.265 1.100 7.150 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.2489 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.710 4.555 1.295 ;
        RECT  3.555 1.205 4.445 1.295 ;
        RECT  3.445 0.710 3.555 1.295 ;
        RECT  2.355 1.205 3.445 1.295 ;
        RECT  2.245 0.710 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.125 -0.165 10.200 0.165 ;
        RECT  10.015 -0.165 10.125 0.690 ;
        RECT  0.000 -0.165 10.015 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.125 1.635 10.200 1.965 ;
        RECT  10.015 1.110 10.125 1.965 ;
        RECT  3.175 1.635 10.015 1.965 ;
        RECT  2.985 1.390 3.175 1.965 ;
        RECT  1.435 1.635 2.985 1.965 ;
        RECT  1.245 1.445 1.435 1.965 ;
        RECT  0.185 1.635 1.245 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.750 0.325 9.905 0.690 ;
        RECT  7.750 1.100 9.905 1.475 ;
        RECT  5.265 0.325 7.050 0.695 ;
        RECT  5.265 1.100 7.050 1.475 ;
        RECT  7.960 0.800 9.970 0.940 ;
        RECT  5.175 0.805 6.990 0.945 ;
        RECT  5.035 0.300 5.175 1.525 ;
        RECT  3.215 0.300 5.035 0.440 ;
        RECT  3.455 1.385 5.035 1.525 ;
        RECT  4.845 0.530 4.945 0.895 ;
        RECT  4.050 0.530 4.845 0.620 ;
        RECT  3.950 0.530 4.050 0.895 ;
        RECT  3.250 0.530 3.950 0.620 ;
        RECT  3.150 0.530 3.250 1.115 ;
        RECT  2.860 1.015 3.150 1.115 ;
        RECT  2.760 0.475 2.860 1.115 ;
        RECT  2.720 1.015 2.760 1.115 ;
        RECT  2.550 0.275 2.650 0.895 ;
        RECT  1.670 0.275 2.550 0.365 ;
        RECT  2.090 1.390 2.440 1.490 ;
        RECT  2.090 0.505 2.430 0.615 ;
        RECT  2.000 0.505 2.090 1.490 ;
        RECT  1.940 0.835 2.000 1.025 ;
        RECT  1.850 0.505 1.890 0.705 ;
        RECT  1.850 1.265 1.890 1.515 ;
        RECT  1.790 0.505 1.850 1.515 ;
        RECT  1.760 0.505 1.790 1.355 ;
        RECT  1.135 1.265 1.760 1.355 ;
        RECT  1.580 0.275 1.670 1.155 ;
        RECT  1.485 0.275 1.580 0.450 ;
        RECT  1.270 1.055 1.580 1.155 ;
        RECT  1.370 0.545 1.470 0.785 ;
        RECT  1.070 0.545 1.370 0.635 ;
        RECT  1.170 0.905 1.270 1.155 ;
        RECT  1.040 1.265 1.135 1.495 ;
        RECT  0.970 0.310 1.070 1.155 ;
        RECT  0.730 1.385 1.040 1.495 ;
        RECT  0.805 0.310 0.970 0.420 ;
        RECT  0.930 1.055 0.970 1.155 ;
        RECT  0.820 1.055 0.930 1.295 ;
        RECT  0.730 0.535 0.880 0.645 ;
        RECT  0.640 0.535 0.730 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD20

MACRO CKLHQD24
    CLASS CORE ;
    FOREIGN CKLHQD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 2.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.650 0.325 11.505 0.690 ;
        RECT  8.650 1.100 11.505 1.475 ;
        RECT  8.150 0.325 8.650 1.475 ;
        RECT  5.865 0.325 8.150 0.695 ;
        RECT  5.865 1.100 8.150 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.2955 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.445 0.710 5.545 1.295 ;
        RECT  4.555 1.205 5.445 1.295 ;
        RECT  4.445 0.710 4.555 1.295 ;
        RECT  3.555 1.205 4.445 1.295 ;
        RECT  3.445 0.710 3.555 1.295 ;
        RECT  2.355 1.205 3.445 1.295 ;
        RECT  2.245 0.710 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.725 -0.165 11.800 0.165 ;
        RECT  11.615 -0.165 11.725 0.690 ;
        RECT  0.000 -0.165 11.615 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.725 1.635 11.800 1.965 ;
        RECT  11.615 1.110 11.725 1.965 ;
        RECT  3.175 1.635 11.615 1.965 ;
        RECT  2.985 1.390 3.175 1.965 ;
        RECT  1.435 1.635 2.985 1.965 ;
        RECT  1.245 1.445 1.435 1.965 ;
        RECT  0.185 1.635 1.245 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.750 0.325 11.505 0.690 ;
        RECT  8.750 1.100 11.505 1.475 ;
        RECT  5.865 0.325 8.050 0.695 ;
        RECT  5.865 1.100 8.050 1.475 ;
        RECT  8.920 0.800 11.330 0.940 ;
        RECT  5.775 0.805 7.980 0.945 ;
        RECT  5.760 0.310 5.775 0.945 ;
        RECT  5.635 0.310 5.760 1.495 ;
        RECT  3.215 0.310 5.635 0.420 ;
        RECT  3.455 1.385 5.635 1.495 ;
        RECT  4.845 0.530 4.955 0.895 ;
        RECT  4.050 0.530 4.845 0.620 ;
        RECT  3.950 0.530 4.050 0.895 ;
        RECT  3.250 0.530 3.950 0.620 ;
        RECT  3.150 0.530 3.250 1.115 ;
        RECT  2.860 1.015 3.150 1.115 ;
        RECT  2.760 0.475 2.860 1.115 ;
        RECT  2.720 1.015 2.760 1.115 ;
        RECT  2.550 0.275 2.650 0.915 ;
        RECT  1.670 0.275 2.550 0.365 ;
        RECT  2.090 1.390 2.440 1.490 ;
        RECT  2.090 0.505 2.430 0.615 ;
        RECT  2.000 0.505 2.090 1.490 ;
        RECT  1.940 0.835 2.000 1.025 ;
        RECT  1.850 0.505 1.890 0.705 ;
        RECT  1.850 1.265 1.890 1.515 ;
        RECT  1.790 0.505 1.850 1.515 ;
        RECT  1.760 0.505 1.790 1.355 ;
        RECT  1.135 1.265 1.760 1.355 ;
        RECT  1.580 0.275 1.670 1.155 ;
        RECT  1.485 0.275 1.580 0.450 ;
        RECT  1.270 1.055 1.580 1.155 ;
        RECT  1.370 0.545 1.470 0.785 ;
        RECT  1.070 0.545 1.370 0.635 ;
        RECT  1.170 0.905 1.270 1.155 ;
        RECT  1.040 1.265 1.135 1.495 ;
        RECT  0.970 0.310 1.070 1.155 ;
        RECT  0.730 1.385 1.040 1.495 ;
        RECT  0.805 0.310 0.970 0.420 ;
        RECT  0.930 1.055 0.970 1.155 ;
        RECT  0.820 1.055 0.930 1.295 ;
        RECT  0.730 0.535 0.880 0.645 ;
        RECT  0.640 0.535 0.730 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD24

MACRO CKLHQD3
    CLASS CORE ;
    FOREIGN CKLHQD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.3270 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.310 4.350 0.690 ;
        RECT  4.250 1.110 4.350 1.490 ;
        RECT  3.950 0.310 4.250 1.490 ;
        RECT  3.715 0.310 3.950 0.690 ;
        RECT  3.715 1.110 3.950 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0739 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.710 3.350 1.295 ;
        RECT  2.355 1.205 3.250 1.295 ;
        RECT  2.245 0.745 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.540 -0.165 4.400 0.165 ;
        RECT  3.350 -0.165 3.540 0.415 ;
        RECT  0.000 -0.165 3.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.475 1.635 4.400 1.965 ;
        RECT  1.265 1.445 1.475 1.965 ;
        RECT  0.185 1.635 1.265 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.715 0.310 3.850 0.690 ;
        RECT  3.715 1.110 3.850 1.490 ;
        RECT  3.500 0.505 3.600 1.490 ;
        RECT  3.025 0.505 3.500 0.615 ;
        RECT  3.185 1.390 3.500 1.490 ;
        RECT  2.960 0.725 3.050 1.115 ;
        RECT  2.590 1.025 2.960 1.115 ;
        RECT  2.780 0.275 2.870 0.905 ;
        RECT  1.700 0.275 2.780 0.365 ;
        RECT  2.700 0.735 2.780 0.905 ;
        RECT  2.590 0.475 2.670 0.645 ;
        RECT  2.500 0.475 2.590 1.115 ;
        RECT  2.120 1.390 2.470 1.490 ;
        RECT  2.120 0.475 2.410 0.645 ;
        RECT  2.030 0.475 2.120 1.490 ;
        RECT  1.970 0.835 2.030 1.025 ;
        RECT  1.880 0.505 1.920 0.705 ;
        RECT  1.880 1.265 1.920 1.515 ;
        RECT  1.820 0.505 1.880 1.515 ;
        RECT  1.790 0.505 1.820 1.355 ;
        RECT  1.150 1.265 1.790 1.355 ;
        RECT  1.610 0.275 1.700 1.155 ;
        RECT  1.525 0.275 1.610 0.450 ;
        RECT  1.295 1.055 1.610 1.155 ;
        RECT  1.400 0.545 1.500 0.785 ;
        RECT  1.070 0.545 1.400 0.635 ;
        RECT  1.195 0.885 1.295 1.155 ;
        RECT  1.050 1.265 1.150 1.495 ;
        RECT  0.970 0.315 1.070 1.155 ;
        RECT  0.740 1.385 1.050 1.495 ;
        RECT  0.805 0.315 0.970 0.425 ;
        RECT  0.940 1.055 0.970 1.155 ;
        RECT  0.830 1.055 0.940 1.295 ;
        RECT  0.740 0.555 0.880 0.665 ;
        RECT  0.640 0.555 0.740 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD3

MACRO CKLHQD4
    CLASS CORE ;
    FOREIGN CKLHQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.310 4.750 0.690 ;
        RECT  4.650 1.110 4.750 1.490 ;
        RECT  4.350 0.310 4.650 1.490 ;
        RECT  4.065 0.310 4.350 0.690 ;
        RECT  4.065 1.110 4.350 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.1381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.710 3.355 1.295 ;
        RECT  2.355 1.205 3.245 1.295 ;
        RECT  2.245 0.745 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 1.635 5.000 1.965 ;
        RECT  3.760 1.390 3.950 1.965 ;
        RECT  2.945 1.635 3.760 1.965 ;
        RECT  2.755 1.390 2.945 1.965 ;
        RECT  1.475 1.635 2.755 1.965 ;
        RECT  1.265 1.445 1.475 1.965 ;
        RECT  0.185 1.635 1.265 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.065 0.310 4.250 0.690 ;
        RECT  4.065 1.110 4.250 1.490 ;
        RECT  3.950 0.800 4.100 0.900 ;
        RECT  3.850 0.310 3.950 1.295 ;
        RECT  3.025 0.310 3.850 0.420 ;
        RECT  3.555 1.205 3.850 1.295 ;
        RECT  3.660 0.530 3.750 0.940 ;
        RECT  3.050 0.530 3.660 0.620 ;
        RECT  3.445 1.205 3.555 1.490 ;
        RECT  3.255 1.390 3.445 1.490 ;
        RECT  2.960 0.530 3.050 1.115 ;
        RECT  2.590 1.025 2.960 1.115 ;
        RECT  2.780 0.275 2.870 0.905 ;
        RECT  1.700 0.275 2.780 0.365 ;
        RECT  2.700 0.735 2.780 0.905 ;
        RECT  2.590 0.475 2.670 0.645 ;
        RECT  2.500 0.475 2.590 1.115 ;
        RECT  2.120 1.390 2.470 1.490 ;
        RECT  2.120 0.475 2.410 0.645 ;
        RECT  2.030 0.475 2.120 1.490 ;
        RECT  1.970 0.835 2.030 1.025 ;
        RECT  1.880 0.505 1.920 0.705 ;
        RECT  1.880 1.265 1.920 1.515 ;
        RECT  1.820 0.505 1.880 1.515 ;
        RECT  1.790 0.505 1.820 1.355 ;
        RECT  1.150 1.265 1.790 1.355 ;
        RECT  1.610 0.275 1.700 1.155 ;
        RECT  1.525 0.275 1.610 0.450 ;
        RECT  1.295 1.055 1.610 1.155 ;
        RECT  1.400 0.545 1.500 0.785 ;
        RECT  1.070 0.545 1.400 0.635 ;
        RECT  1.195 0.885 1.295 1.155 ;
        RECT  1.050 1.265 1.150 1.495 ;
        RECT  0.970 0.315 1.070 1.155 ;
        RECT  0.740 1.385 1.050 1.495 ;
        RECT  0.805 0.315 0.970 0.425 ;
        RECT  0.940 1.055 0.970 1.155 ;
        RECT  0.830 1.055 0.940 1.295 ;
        RECT  0.740 0.555 0.880 0.665 ;
        RECT  0.640 0.555 0.740 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD4

MACRO CKLHQD6
    CLASS CORE ;
    FOREIGN CKLHQD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.5460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.310 5.215 0.690 ;
        RECT  4.850 1.110 5.215 1.490 ;
        RECT  4.550 0.310 4.850 1.490 ;
        RECT  4.065 0.310 4.550 0.690 ;
        RECT  4.065 1.110 4.550 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.1381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.710 3.355 1.295 ;
        RECT  2.355 1.205 3.245 1.295 ;
        RECT  2.245 0.745 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.435 -0.165 5.600 0.165 ;
        RECT  5.325 -0.165 5.435 0.690 ;
        RECT  0.000 -0.165 5.325 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.435 1.635 5.600 1.965 ;
        RECT  5.325 1.110 5.435 1.965 ;
        RECT  3.950 1.635 5.325 1.965 ;
        RECT  3.760 1.390 3.950 1.965 ;
        RECT  2.945 1.635 3.760 1.965 ;
        RECT  2.755 1.390 2.945 1.965 ;
        RECT  1.475 1.635 2.755 1.965 ;
        RECT  1.265 1.445 1.475 1.965 ;
        RECT  0.185 1.635 1.265 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.950 0.310 5.215 0.690 ;
        RECT  4.950 1.110 5.215 1.490 ;
        RECT  4.065 0.310 4.450 0.690 ;
        RECT  4.065 1.110 4.450 1.490 ;
        RECT  3.950 0.800 4.100 0.900 ;
        RECT  3.850 0.310 3.950 1.295 ;
        RECT  3.015 0.310 3.850 0.420 ;
        RECT  3.555 1.205 3.850 1.295 ;
        RECT  3.660 0.530 3.750 0.940 ;
        RECT  3.050 0.530 3.660 0.620 ;
        RECT  3.445 1.205 3.555 1.490 ;
        RECT  3.255 1.390 3.445 1.490 ;
        RECT  2.960 0.530 3.050 1.115 ;
        RECT  2.590 1.025 2.960 1.115 ;
        RECT  2.780 0.275 2.870 0.905 ;
        RECT  1.700 0.275 2.780 0.365 ;
        RECT  2.700 0.735 2.780 0.905 ;
        RECT  2.590 0.475 2.670 0.645 ;
        RECT  2.500 0.475 2.590 1.115 ;
        RECT  2.120 1.390 2.470 1.490 ;
        RECT  2.120 0.475 2.410 0.645 ;
        RECT  2.030 0.475 2.120 1.490 ;
        RECT  1.970 0.835 2.030 1.025 ;
        RECT  1.880 0.505 1.920 0.705 ;
        RECT  1.880 1.265 1.920 1.515 ;
        RECT  1.820 0.505 1.880 1.515 ;
        RECT  1.790 0.505 1.820 1.355 ;
        RECT  1.150 1.265 1.790 1.355 ;
        RECT  1.610 0.275 1.700 1.155 ;
        RECT  1.525 0.275 1.610 0.450 ;
        RECT  1.295 1.055 1.610 1.155 ;
        RECT  1.400 0.545 1.500 0.785 ;
        RECT  1.070 0.545 1.400 0.635 ;
        RECT  1.195 0.885 1.295 1.155 ;
        RECT  1.050 1.265 1.150 1.495 ;
        RECT  0.970 0.315 1.070 1.155 ;
        RECT  0.740 1.385 1.050 1.495 ;
        RECT  0.805 0.315 0.970 0.425 ;
        RECT  0.940 1.055 0.970 1.155 ;
        RECT  0.830 1.055 0.940 1.295 ;
        RECT  0.740 0.555 0.880 0.665 ;
        RECT  0.640 0.555 0.740 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD6

MACRO CKLHQD8
    CLASS CORE ;
    FOREIGN CKLHQD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.955 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.325 5.715 0.695 ;
        RECT  5.050 1.105 5.715 1.475 ;
        RECT  4.550 0.325 5.050 1.475 ;
        RECT  4.065 0.325 4.550 0.695 ;
        RECT  4.065 1.105 4.550 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 1.090 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.1381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.710 3.355 1.295 ;
        RECT  2.355 1.205 3.245 1.295 ;
        RECT  2.245 0.745 2.355 1.295 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 6.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 1.635 6.000 1.965 ;
        RECT  3.760 1.390 3.950 1.965 ;
        RECT  2.945 1.635 3.760 1.965 ;
        RECT  2.755 1.390 2.945 1.965 ;
        RECT  1.475 1.635 2.755 1.965 ;
        RECT  1.265 1.445 1.475 1.965 ;
        RECT  0.185 1.635 1.265 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.150 0.325 5.715 0.695 ;
        RECT  5.150 1.105 5.715 1.475 ;
        RECT  4.065 0.325 4.450 0.695 ;
        RECT  4.065 1.105 4.450 1.475 ;
        RECT  5.250 0.805 5.680 0.940 ;
        RECT  3.975 0.805 4.385 0.940 ;
        RECT  3.830 0.300 3.975 1.295 ;
        RECT  3.025 0.300 3.830 0.440 ;
        RECT  3.645 1.170 3.830 1.295 ;
        RECT  3.630 0.530 3.740 0.940 ;
        RECT  3.535 1.170 3.645 1.520 ;
        RECT  3.050 0.530 3.630 0.620 ;
        RECT  3.255 1.390 3.535 1.520 ;
        RECT  2.960 0.530 3.050 1.115 ;
        RECT  2.590 1.025 2.960 1.115 ;
        RECT  2.780 0.275 2.870 0.905 ;
        RECT  1.700 0.275 2.780 0.365 ;
        RECT  2.700 0.735 2.780 0.905 ;
        RECT  2.590 0.475 2.670 0.645 ;
        RECT  2.500 0.475 2.590 1.115 ;
        RECT  2.120 1.390 2.470 1.490 ;
        RECT  2.120 0.475 2.410 0.645 ;
        RECT  2.030 0.475 2.120 1.490 ;
        RECT  1.970 0.835 2.030 1.025 ;
        RECT  1.880 0.505 1.920 0.705 ;
        RECT  1.880 1.265 1.920 1.515 ;
        RECT  1.820 0.505 1.880 1.515 ;
        RECT  1.790 0.505 1.820 1.355 ;
        RECT  1.150 1.265 1.790 1.355 ;
        RECT  1.610 0.275 1.700 1.155 ;
        RECT  1.525 0.275 1.610 0.450 ;
        RECT  1.295 1.055 1.610 1.155 ;
        RECT  1.400 0.545 1.500 0.785 ;
        RECT  1.070 0.545 1.400 0.635 ;
        RECT  1.195 0.885 1.295 1.155 ;
        RECT  1.050 1.265 1.150 1.495 ;
        RECT  0.970 0.315 1.070 1.155 ;
        RECT  0.740 1.385 1.050 1.495 ;
        RECT  0.805 0.315 0.970 0.425 ;
        RECT  0.940 1.055 0.970 1.155 ;
        RECT  0.830 1.055 0.940 1.295 ;
        RECT  0.740 0.555 0.880 0.665 ;
        RECT  0.640 0.555 0.740 1.495 ;
        RECT  0.185 0.310 0.715 0.420 ;
        RECT  0.075 0.310 0.185 0.565 ;
    END
END CKLHQD8

MACRO CKLNQD1
    CLASS CORE ;
    FOREIGN CKLNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.1170 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.465 3.550 1.490 ;
        RECT  3.415 0.465 3.450 0.675 ;
        RECT  3.415 1.040 3.450 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0622 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.900 2.555 1.300 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 3.600 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.575 1.635 3.600 1.965 ;
        RECT  1.365 1.445 1.575 1.965 ;
        RECT  0.190 1.635 1.365 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.305 0.760 3.360 0.950 ;
        RECT  3.215 0.760 3.305 1.445 ;
        RECT  2.825 1.335 3.215 1.445 ;
        RECT  3.010 0.275 3.120 1.135 ;
        RECT  1.810 0.275 3.010 0.365 ;
        RECT  2.715 0.455 2.825 1.445 ;
        RECT  2.300 0.505 2.605 0.615 ;
        RECT  2.300 1.390 2.580 1.490 ;
        RECT  2.210 0.505 2.300 1.490 ;
        RECT  2.105 0.750 2.210 0.920 ;
        RECT  2.015 0.465 2.045 0.655 ;
        RECT  2.015 1.265 2.030 1.520 ;
        RECT  1.920 0.465 2.015 1.520 ;
        RECT  1.140 1.265 1.920 1.355 ;
        RECT  1.710 0.275 1.810 1.175 ;
        RECT  1.675 0.275 1.710 0.485 ;
        RECT  1.360 1.060 1.710 1.175 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.815 1.360 1.175 ;
        RECT  1.140 0.595 1.250 0.705 ;
        RECT  1.050 0.595 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD1

MACRO CKLNQD12
    CLASS CORE ;
    FOREIGN CKLNQD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.8880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.325 6.515 0.690 ;
        RECT  5.450 1.100 6.515 1.475 ;
        RECT  4.950 0.325 5.450 1.475 ;
        RECT  3.875 0.325 4.950 0.690 ;
        RECT  3.875 1.100 4.950 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0974 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.565 1.135 ;
        RECT  2.555 1.025 3.450 1.135 ;
        RECT  2.445 0.700 2.555 1.135 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 -0.165 6.800 0.165 ;
        RECT  3.550 -0.165 3.720 0.390 ;
        RECT  0.520 -0.165 3.550 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.635 6.800 1.965 ;
        RECT  1.330 1.445 1.540 1.965 ;
        RECT  0.190 1.635 1.330 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.550 0.325 6.515 0.690 ;
        RECT  5.550 1.100 6.515 1.475 ;
        RECT  3.875 0.325 4.850 0.690 ;
        RECT  3.875 1.100 4.850 1.475 ;
        RECT  5.590 0.800 6.520 0.940 ;
        RECT  3.785 0.800 4.785 0.940 ;
        RECT  3.655 0.480 3.785 1.420 ;
        RECT  3.055 0.480 3.655 0.620 ;
        RECT  2.815 1.280 3.655 1.420 ;
        RECT  2.940 0.780 3.250 0.890 ;
        RECT  2.830 0.275 2.940 0.890 ;
        RECT  1.810 0.275 2.830 0.365 ;
        RECT  2.300 0.500 2.585 0.610 ;
        RECT  2.300 1.310 2.550 1.420 ;
        RECT  2.210 0.500 2.300 1.420 ;
        RECT  2.100 0.750 2.210 0.920 ;
        RECT  2.010 0.465 2.045 0.655 ;
        RECT  1.920 0.465 2.010 1.520 ;
        RECT  1.890 1.265 1.920 1.520 ;
        RECT  1.140 1.265 1.890 1.355 ;
        RECT  1.710 0.275 1.810 1.175 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.060 1.710 1.175 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.785 1.360 1.175 ;
        RECT  1.140 0.565 1.250 0.675 ;
        RECT  1.050 0.565 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD12

MACRO CKLNQD16
    CLASS CORE ;
    FOREIGN CKLNQD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.325 8.105 0.690 ;
        RECT  6.650 1.100 8.105 1.475 ;
        RECT  6.150 0.325 6.650 1.475 ;
        RECT  4.445 0.325 6.150 0.690 ;
        RECT  4.445 1.100 6.150 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.1321 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.005 0.750 4.115 1.090 ;
        RECT  2.555 0.910 4.005 1.090 ;
        RECT  2.445 0.910 2.555 1.300 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 8.400 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.575 1.635 8.400 1.965 ;
        RECT  1.365 1.445 1.575 1.965 ;
        RECT  0.190 1.635 1.365 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.750 0.325 8.105 0.690 ;
        RECT  6.750 1.100 8.105 1.475 ;
        RECT  4.445 0.325 6.050 0.690 ;
        RECT  4.445 1.100 6.050 1.475 ;
        RECT  6.810 0.800 8.220 0.940 ;
        RECT  4.355 0.800 5.980 0.940 ;
        RECT  4.205 0.485 4.355 1.410 ;
        RECT  2.660 0.485 4.205 0.625 ;
        RECT  2.845 1.270 4.205 1.410 ;
        RECT  2.730 0.275 3.815 0.390 ;
        RECT  1.810 0.275 2.730 0.365 ;
        RECT  2.300 1.390 2.580 1.495 ;
        RECT  2.445 0.455 2.555 0.655 ;
        RECT  2.300 0.545 2.445 0.655 ;
        RECT  2.210 0.545 2.300 1.495 ;
        RECT  2.100 0.750 2.210 0.920 ;
        RECT  2.010 0.465 2.045 0.655 ;
        RECT  2.010 1.265 2.030 1.520 ;
        RECT  1.920 0.465 2.010 1.520 ;
        RECT  1.140 1.265 1.920 1.355 ;
        RECT  1.710 0.275 1.810 1.175 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.060 1.710 1.175 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.815 1.360 1.175 ;
        RECT  1.140 0.595 1.250 0.705 ;
        RECT  1.050 0.595 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD16

MACRO CKLNQD2
    CLASS CORE ;
    FOREIGN CKLNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.090 ;
        RECT  0.180 0.710 0.245 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.1480 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.460 0.510 3.555 1.140 ;
        RECT  3.445 0.510 3.460 1.490 ;
        RECT  3.310 0.510 3.445 0.620 ;
        RECT  3.350 1.040 3.445 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.615 0.640 0.725 ;
        RECT  0.445 0.615 0.555 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0626 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.700 2.550 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 3.800 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 1.635 3.800 1.965 ;
        RECT  3.610 1.250 3.720 1.965 ;
        RECT  1.490 1.635 3.610 1.965 ;
        RECT  1.280 1.445 1.490 1.965 ;
        RECT  0.190 1.635 1.280 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.255 0.760 3.335 0.930 ;
        RECT  3.165 0.760 3.255 1.355 ;
        RECT  2.770 1.245 3.165 1.355 ;
        RECT  2.945 0.275 3.050 1.135 ;
        RECT  1.805 0.275 2.945 0.365 ;
        RECT  2.660 0.455 2.770 1.355 ;
        RECT  2.240 0.455 2.550 0.565 ;
        RECT  2.240 1.270 2.495 1.370 ;
        RECT  2.150 0.455 2.240 1.370 ;
        RECT  2.075 0.910 2.150 1.080 ;
        RECT  1.985 0.510 2.005 0.700 ;
        RECT  1.895 0.510 1.985 1.520 ;
        RECT  1.860 1.265 1.895 1.520 ;
        RECT  1.140 1.265 1.860 1.355 ;
        RECT  1.710 0.275 1.805 1.175 ;
        RECT  1.360 1.065 1.710 1.175 ;
        RECT  1.520 0.330 1.620 0.940 ;
        RECT  0.960 0.330 1.520 0.440 ;
        RECT  1.250 0.785 1.360 1.175 ;
        RECT  1.140 0.565 1.250 0.675 ;
        RECT  1.050 0.565 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.645 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD2

MACRO CKLNQD20
    CLASS CORE ;
    FOREIGN CKLNQD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.4800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.325 9.515 0.690 ;
        RECT  7.450 1.100 9.515 1.475 ;
        RECT  6.950 0.325 7.450 1.475 ;
        RECT  4.875 0.325 6.950 0.690 ;
        RECT  4.875 1.100 6.950 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.1664 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.735 4.560 1.090 ;
        RECT  2.555 0.955 4.450 1.090 ;
        RECT  2.445 0.900 2.555 1.300 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.490 -0.165 9.800 0.165 ;
        RECT  0.380 -0.165 0.490 0.325 ;
        RECT  0.000 -0.165 0.380 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.635 9.800 1.965 ;
        RECT  1.335 1.445 1.545 1.965 ;
        RECT  0.190 1.635 1.335 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.550 0.325 9.515 0.690 ;
        RECT  7.550 1.100 9.515 1.475 ;
        RECT  4.875 0.325 6.850 0.690 ;
        RECT  4.875 1.100 6.850 1.475 ;
        RECT  7.610 0.800 9.490 0.940 ;
        RECT  4.785 0.800 6.775 0.940 ;
        RECT  4.650 0.485 4.785 1.430 ;
        RECT  3.085 0.485 4.650 0.625 ;
        RECT  2.815 1.290 4.650 1.430 ;
        RECT  2.810 0.755 4.285 0.865 ;
        RECT  2.720 0.275 2.810 0.865 ;
        RECT  1.810 0.275 2.720 0.365 ;
        RECT  2.300 0.505 2.605 0.615 ;
        RECT  2.300 1.390 2.550 1.495 ;
        RECT  2.210 0.505 2.300 1.495 ;
        RECT  2.100 0.750 2.210 0.920 ;
        RECT  2.000 0.465 2.045 0.655 ;
        RECT  1.900 0.465 2.000 1.520 ;
        RECT  1.890 1.265 1.900 1.520 ;
        RECT  1.140 1.265 1.890 1.355 ;
        RECT  1.710 0.275 1.810 1.160 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.050 1.710 1.160 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.785 1.360 1.160 ;
        RECT  1.140 0.565 1.250 0.675 ;
        RECT  1.050 0.565 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD20

MACRO CKLNQD24
    CLASS CORE ;
    FOREIGN CKLNQD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.7760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 0.325 10.515 0.690 ;
        RECT  8.050 1.100 10.515 1.475 ;
        RECT  7.550 0.325 8.050 1.475 ;
        RECT  4.870 0.325 7.550 0.690 ;
        RECT  4.870 1.100 7.550 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.1664 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.435 0.710 4.545 1.090 ;
        RECT  2.555 0.955 4.435 1.090 ;
        RECT  2.445 0.900 2.555 1.300 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 10.800 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.635 10.800 1.965 ;
        RECT  1.330 1.445 1.540 1.965 ;
        RECT  0.190 1.635 1.330 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.150 0.325 10.515 0.690 ;
        RECT  8.150 1.100 10.515 1.475 ;
        RECT  4.870 0.325 7.450 0.690 ;
        RECT  4.870 1.100 7.450 1.475 ;
        RECT  8.210 0.800 10.540 0.940 ;
        RECT  4.780 0.800 7.365 0.940 ;
        RECT  4.635 0.480 4.780 1.410 ;
        RECT  3.065 0.480 4.635 0.620 ;
        RECT  2.810 1.270 4.635 1.410 ;
        RECT  2.840 0.755 4.280 0.865 ;
        RECT  2.750 0.275 2.840 0.865 ;
        RECT  1.810 0.275 2.750 0.365 ;
        RECT  2.300 0.505 2.605 0.615 ;
        RECT  2.300 1.390 2.545 1.495 ;
        RECT  2.210 0.505 2.300 1.495 ;
        RECT  2.100 0.750 2.210 0.920 ;
        RECT  2.010 0.465 2.045 0.655 ;
        RECT  1.920 0.465 2.010 1.520 ;
        RECT  1.885 1.265 1.920 1.520 ;
        RECT  1.140 1.265 1.885 1.355 ;
        RECT  1.710 0.275 1.810 1.150 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.050 1.710 1.150 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.815 1.360 1.150 ;
        RECT  1.140 0.595 1.250 0.705 ;
        RECT  1.050 0.595 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD24

MACRO CKLNQD3
    CLASS CORE ;
    FOREIGN CKLNQD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.2770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.455 4.150 0.625 ;
        RECT  3.990 1.040 4.100 1.490 ;
        RECT  3.850 1.040 3.990 1.210 ;
        RECT  3.580 0.455 3.850 1.210 ;
        RECT  3.550 0.455 3.580 1.490 ;
        RECT  3.420 0.455 3.550 0.625 ;
        RECT  3.450 1.040 3.550 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0621 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.900 2.555 1.300 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.165 4.200 0.165 ;
        RECT  3.195 -0.165 3.310 0.675 ;
        RECT  0.520 -0.165 3.195 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.855 1.635 4.200 1.965 ;
        RECT  3.715 1.320 3.855 1.965 ;
        RECT  3.325 1.635 3.715 1.965 ;
        RECT  3.155 1.505 3.325 1.965 ;
        RECT  1.575 1.635 3.155 1.965 ;
        RECT  1.365 1.445 1.575 1.965 ;
        RECT  0.190 1.635 1.365 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.950 0.455 4.150 0.625 ;
        RECT  3.990 1.040 4.100 1.490 ;
        RECT  3.950 1.040 3.990 1.210 ;
        RECT  3.420 0.455 3.450 0.625 ;
        RECT  3.305 0.790 3.425 0.900 ;
        RECT  3.215 0.790 3.305 1.415 ;
        RECT  2.820 1.305 3.215 1.415 ;
        RECT  2.995 0.275 3.105 1.135 ;
        RECT  1.810 0.275 2.995 0.365 ;
        RECT  2.710 0.465 2.820 1.415 ;
        RECT  2.300 0.515 2.600 0.625 ;
        RECT  2.300 1.390 2.565 1.490 ;
        RECT  2.210 0.515 2.300 1.490 ;
        RECT  2.105 0.750 2.210 0.920 ;
        RECT  2.015 0.465 2.045 0.655 ;
        RECT  2.015 1.265 2.030 1.520 ;
        RECT  1.920 0.465 2.015 1.520 ;
        RECT  1.140 1.265 1.920 1.355 ;
        RECT  1.710 0.275 1.810 1.175 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.060 1.710 1.175 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.815 1.360 1.175 ;
        RECT  1.140 0.595 1.250 0.705 ;
        RECT  1.050 0.595 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD3

MACRO CKLNQD4
    CLASS CORE ;
    FOREIGN CKLNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.2960 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.510 4.070 0.690 ;
        RECT  3.850 1.110 4.070 1.490 ;
        RECT  3.550 0.510 3.850 1.490 ;
        RECT  3.360 0.510 3.550 0.690 ;
        RECT  3.400 1.110 3.550 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0621 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.900 2.555 1.300 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.300 -0.165 4.400 0.165 ;
        RECT  4.190 -0.165 4.300 0.675 ;
        RECT  0.520 -0.165 4.190 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.635 4.400 1.965 ;
        RECT  4.180 1.040 4.290 1.965 ;
        RECT  1.575 1.635 4.180 1.965 ;
        RECT  1.365 1.445 1.575 1.965 ;
        RECT  0.190 1.635 1.365 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.950 0.510 4.070 0.690 ;
        RECT  3.950 1.110 4.070 1.490 ;
        RECT  3.360 0.510 3.450 0.690 ;
        RECT  3.400 1.110 3.450 1.490 ;
        RECT  3.305 0.800 3.420 0.900 ;
        RECT  3.215 0.800 3.305 1.420 ;
        RECT  2.820 1.310 3.215 1.420 ;
        RECT  2.995 0.275 3.105 1.135 ;
        RECT  1.810 0.275 2.995 0.365 ;
        RECT  2.710 0.465 2.820 1.420 ;
        RECT  2.300 0.515 2.600 0.625 ;
        RECT  2.300 1.390 2.565 1.490 ;
        RECT  2.210 0.515 2.300 1.490 ;
        RECT  2.105 0.750 2.210 0.920 ;
        RECT  2.015 0.465 2.045 0.655 ;
        RECT  2.015 1.265 2.030 1.520 ;
        RECT  1.920 0.465 2.015 1.520 ;
        RECT  1.140 1.265 1.920 1.355 ;
        RECT  1.710 0.275 1.810 1.175 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.060 1.710 1.175 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.815 1.360 1.175 ;
        RECT  1.140 0.595 1.250 0.705 ;
        RECT  1.050 0.595 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD4

MACRO CKLNQD6
    CLASS CORE ;
    FOREIGN CKLNQD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.4440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.510 5.070 0.690 ;
        RECT  4.650 1.110 5.070 1.490 ;
        RECT  4.350 0.510 4.650 1.490 ;
        RECT  3.870 0.510 4.350 0.690 ;
        RECT  3.900 1.110 4.350 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0973 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.730 3.600 0.940 ;
        RECT  3.450 0.730 3.550 1.135 ;
        RECT  2.555 1.025 3.450 1.135 ;
        RECT  2.445 0.900 2.555 1.300 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.290 -0.165 5.400 0.165 ;
        RECT  5.180 -0.165 5.290 0.675 ;
        RECT  3.755 -0.165 5.180 0.165 ;
        RECT  3.585 -0.165 3.755 0.405 ;
        RECT  0.520 -0.165 3.585 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.290 1.635 5.400 1.965 ;
        RECT  5.180 1.040 5.290 1.965 ;
        RECT  1.575 1.635 5.180 1.965 ;
        RECT  1.365 1.445 1.575 1.965 ;
        RECT  0.190 1.635 1.365 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.750 0.510 5.070 0.690 ;
        RECT  4.750 1.110 5.070 1.490 ;
        RECT  3.870 0.510 4.250 0.690 ;
        RECT  3.900 1.110 4.250 1.490 ;
        RECT  3.780 0.800 4.245 0.900 ;
        RECT  3.690 0.515 3.780 1.420 ;
        RECT  3.090 0.515 3.690 0.625 ;
        RECT  2.850 1.310 3.690 1.420 ;
        RECT  2.975 0.780 3.285 0.890 ;
        RECT  2.865 0.275 2.975 0.890 ;
        RECT  1.810 0.275 2.865 0.365 ;
        RECT  2.300 0.515 2.600 0.625 ;
        RECT  2.300 1.390 2.565 1.490 ;
        RECT  2.210 0.515 2.300 1.490 ;
        RECT  2.105 0.750 2.210 0.920 ;
        RECT  2.015 0.465 2.045 0.655 ;
        RECT  2.015 1.265 2.030 1.520 ;
        RECT  1.920 0.465 2.015 1.520 ;
        RECT  1.140 1.265 1.920 1.355 ;
        RECT  1.710 0.275 1.810 1.175 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.060 1.710 1.175 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.815 1.360 1.175 ;
        RECT  1.140 0.595 1.250 0.705 ;
        RECT  1.050 0.595 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD6

MACRO CKLNQD8
    CLASS CORE ;
    FOREIGN CKLNQD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.180 0.710 0.250 0.940 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.5920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.325 5.515 0.690 ;
        RECT  4.850 1.100 5.515 1.475 ;
        RECT  4.350 0.325 4.850 1.475 ;
        RECT  3.875 0.325 4.350 0.690 ;
        RECT  3.875 1.100 4.350 1.475 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0457 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.615 0.640 0.725 ;
        RECT  0.450 0.615 0.550 1.090 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0973 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.560 1.135 ;
        RECT  2.555 1.025 3.450 1.135 ;
        RECT  2.445 0.700 2.555 1.135 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.800 0.165 ;
        RECT  0.350 -0.165 0.520 0.325 ;
        RECT  0.000 -0.165 0.350 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.635 5.800 1.965 ;
        RECT  1.330 1.445 1.540 1.965 ;
        RECT  0.190 1.635 1.330 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.950 0.325 5.515 0.690 ;
        RECT  4.950 1.100 5.515 1.475 ;
        RECT  3.875 0.325 4.250 0.690 ;
        RECT  3.875 1.100 4.250 1.475 ;
        RECT  5.035 0.800 5.500 0.940 ;
        RECT  3.785 0.800 4.190 0.940 ;
        RECT  3.650 0.480 3.785 1.440 ;
        RECT  3.065 0.480 3.650 0.620 ;
        RECT  2.815 1.295 3.650 1.440 ;
        RECT  2.940 0.780 3.250 0.890 ;
        RECT  2.830 0.275 2.940 0.890 ;
        RECT  1.810 0.275 2.830 0.365 ;
        RECT  2.300 0.480 2.600 0.590 ;
        RECT  2.300 1.310 2.550 1.420 ;
        RECT  2.210 0.480 2.300 1.420 ;
        RECT  2.105 0.750 2.210 0.920 ;
        RECT  1.995 0.465 2.045 0.655 ;
        RECT  1.900 0.465 1.995 1.520 ;
        RECT  1.885 1.265 1.900 1.520 ;
        RECT  1.140 1.265 1.885 1.355 ;
        RECT  1.710 0.275 1.810 1.165 ;
        RECT  1.675 0.275 1.710 0.490 ;
        RECT  1.360 1.050 1.710 1.165 ;
        RECT  1.550 0.625 1.620 0.940 ;
        RECT  1.520 0.330 1.550 0.940 ;
        RECT  1.450 0.330 1.520 0.725 ;
        RECT  0.960 0.330 1.450 0.440 ;
        RECT  1.250 0.785 1.360 1.165 ;
        RECT  1.140 0.565 1.250 0.675 ;
        RECT  1.050 0.565 1.140 1.445 ;
        RECT  0.740 1.355 1.050 1.445 ;
        RECT  0.870 0.330 0.960 1.245 ;
        RECT  0.830 1.035 0.870 1.245 ;
        RECT  0.665 0.315 0.775 0.525 ;
        RECT  0.640 0.835 0.740 1.445 ;
        RECT  0.050 0.415 0.665 0.525 ;
    END
END CKLNQD8

MACRO CKMUX2D0
    CLASS CORE ;
    FOREIGN CKMUX2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.310 1.950 1.490 ;
        RECT  1.825 0.310 1.850 0.600 ;
        RECT  1.815 1.025 1.850 1.490 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0502 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.355 1.100 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0256 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.365 0.700 1.450 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0250 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.630 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.505 -0.165 2.000 0.165 ;
        RECT  0.335 -0.165 0.505 0.575 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.635 2.000 1.965 ;
        RECT  1.515 1.210 1.645 1.965 ;
        RECT  0.515 1.635 1.515 1.965 ;
        RECT  0.345 1.425 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.735 0.730 1.760 0.940 ;
        RECT  1.640 0.275 1.735 0.940 ;
        RECT  1.020 0.275 1.640 0.365 ;
        RECT  1.270 0.455 1.405 0.565 ;
        RECT  1.270 1.190 1.395 1.300 ;
        RECT  1.180 0.455 1.270 1.300 ;
        RECT  0.815 1.425 1.235 1.525 ;
        RECT  1.020 1.020 1.080 1.335 ;
        RECT  0.970 0.275 1.020 1.335 ;
        RECT  0.910 0.275 0.970 1.130 ;
        RECT  0.720 0.465 0.820 1.130 ;
        RECT  0.725 1.240 0.815 1.525 ;
        RECT  0.185 1.240 0.725 1.335 ;
        RECT  0.600 0.465 0.720 0.575 ;
        RECT  0.640 1.030 0.720 1.130 ;
        RECT  0.160 0.425 0.185 0.615 ;
        RECT  0.160 1.240 0.185 1.490 ;
        RECT  0.060 0.425 0.160 1.490 ;
    END
END CKMUX2D0

MACRO CKMUX2D1
    CLASS CORE ;
    FOREIGN CKMUX2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.310 1.950 1.490 ;
        RECT  1.825 0.310 1.850 0.520 ;
        RECT  1.815 1.025 1.850 1.490 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.355 1.100 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.365 0.700 1.450 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.630 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.505 -0.165 2.000 0.165 ;
        RECT  0.335 -0.165 0.505 0.575 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.635 2.000 1.965 ;
        RECT  1.515 1.220 1.650 1.965 ;
        RECT  0.515 1.635 1.515 1.965 ;
        RECT  0.345 1.425 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.735 0.730 1.760 0.940 ;
        RECT  1.640 0.275 1.735 0.940 ;
        RECT  1.020 0.275 1.640 0.365 ;
        RECT  1.270 0.455 1.405 0.565 ;
        RECT  1.270 1.190 1.395 1.300 ;
        RECT  1.180 0.455 1.270 1.300 ;
        RECT  0.815 1.425 1.235 1.525 ;
        RECT  1.020 1.020 1.080 1.335 ;
        RECT  0.970 0.275 1.020 1.335 ;
        RECT  0.910 0.275 0.970 1.130 ;
        RECT  0.720 0.465 0.820 1.130 ;
        RECT  0.725 1.240 0.815 1.525 ;
        RECT  0.185 1.240 0.725 1.335 ;
        RECT  0.600 0.465 0.720 0.575 ;
        RECT  0.640 1.030 0.720 1.130 ;
        RECT  0.160 0.425 0.185 0.615 ;
        RECT  0.160 1.240 0.185 1.490 ;
        RECT  0.060 0.425 0.160 1.490 ;
    END
END CKMUX2D1

MACRO CKMUX2D2
    CLASS CORE ;
    FOREIGN CKMUX2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.305 2.150 1.135 ;
        RECT  1.715 0.305 2.050 0.410 ;
        RECT  1.950 1.035 2.050 1.135 ;
        RECT  1.760 1.035 1.950 1.490 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.355 1.100 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.365 0.700 1.450 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.630 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.505 -0.165 2.200 0.165 ;
        RECT  0.335 -0.165 0.505 0.575 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.635 2.200 1.965 ;
        RECT  1.505 1.255 1.615 1.965 ;
        RECT  0.515 1.635 1.505 1.965 ;
        RECT  0.345 1.425 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.765 0.500 1.875 0.930 ;
        RECT  1.605 0.500 1.765 0.590 ;
        RECT  1.515 0.275 1.605 0.590 ;
        RECT  1.020 0.275 1.515 0.365 ;
        RECT  1.270 0.455 1.405 0.565 ;
        RECT  1.270 1.190 1.395 1.300 ;
        RECT  1.180 0.455 1.270 1.300 ;
        RECT  0.815 1.425 1.235 1.525 ;
        RECT  1.020 1.020 1.080 1.335 ;
        RECT  0.970 0.275 1.020 1.335 ;
        RECT  0.910 0.275 0.970 1.130 ;
        RECT  0.720 0.465 0.820 1.130 ;
        RECT  0.725 1.240 0.815 1.525 ;
        RECT  0.185 1.240 0.725 1.335 ;
        RECT  0.600 0.465 0.720 0.575 ;
        RECT  0.640 1.030 0.720 1.130 ;
        RECT  0.160 0.425 0.185 0.615 ;
        RECT  0.160 1.240 0.185 1.490 ;
        RECT  0.060 0.425 0.160 1.490 ;
    END
END CKMUX2D2

MACRO CKMUX2D4
    CLASS CORE ;
    FOREIGN CKMUX2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.060 0.690 ;
        RECT  3.050 1.030 3.060 1.480 ;
        RECT  2.950 0.275 3.050 1.480 ;
        RECT  2.750 0.595 2.950 1.130 ;
        RECT  2.540 0.595 2.750 0.690 ;
        RECT  2.540 1.030 2.750 1.130 ;
        RECT  2.440 0.275 2.540 0.690 ;
        RECT  2.430 1.030 2.540 1.480 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0557 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.750 1.100 ;
        RECT  1.545 0.755 1.650 0.925 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.700 2.150 1.100 ;
        RECT  2.020 0.700 2.050 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.550 0.900 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.320 -0.165 3.400 0.165 ;
        RECT  3.210 -0.165 3.320 0.705 ;
        RECT  2.800 -0.165 3.210 0.165 ;
        RECT  2.690 -0.165 2.800 0.485 ;
        RECT  0.000 -0.165 2.690 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.635 3.400 1.965 ;
        RECT  3.210 1.030 3.320 1.965 ;
        RECT  2.800 1.635 3.210 1.965 ;
        RECT  2.690 1.285 2.800 1.965 ;
        RECT  2.265 1.635 2.690 1.965 ;
        RECT  2.155 1.285 2.265 1.965 ;
        RECT  0.000 1.635 2.155 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.540 0.595 2.650 0.690 ;
        RECT  2.540 1.030 2.650 1.130 ;
        RECT  2.440 0.275 2.540 0.690 ;
        RECT  2.430 1.030 2.540 1.480 ;
        RECT  2.330 0.780 2.525 0.890 ;
        RECT  2.240 0.275 2.330 0.890 ;
        RECT  0.945 0.275 2.240 0.365 ;
        RECT  1.930 0.500 2.070 0.610 ;
        RECT  1.930 1.295 2.045 1.405 ;
        RECT  1.840 0.500 1.930 1.405 ;
        RECT  1.205 1.315 1.840 1.405 ;
        RECT  1.450 0.475 1.490 0.675 ;
        RECT  1.450 1.015 1.480 1.225 ;
        RECT  1.360 0.475 1.450 1.225 ;
        RECT  1.295 0.755 1.360 0.925 ;
        RECT  1.205 0.455 1.230 0.645 ;
        RECT  1.095 0.455 1.205 1.405 ;
        RECT  0.835 0.275 0.945 1.330 ;
        RECT  0.185 1.170 0.735 1.280 ;
        RECT  0.575 0.280 0.685 0.490 ;
        RECT  0.185 0.400 0.575 0.490 ;
        RECT  0.145 0.280 0.185 0.490 ;
        RECT  0.145 1.055 0.185 1.485 ;
        RECT  0.055 0.280 0.145 1.485 ;
    END
END CKMUX2D4

MACRO CKND0
    CLASS CORE ;
    FOREIGN CKND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.580 0.550 1.110 ;
        RECT  0.425 0.275 0.455 1.490 ;
        RECT  0.345 0.275 0.425 0.695 ;
        RECT  0.345 1.000 0.425 1.490 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0250 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.185 0.930 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 1.635 0.600 1.965 ;
        RECT  0.085 1.220 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END CKND0

MACRO CKND1
    CLASS CORE ;
    FOREIGN CKND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.580 0.550 1.110 ;
        RECT  0.425 0.275 0.455 1.490 ;
        RECT  0.345 0.275 0.425 0.695 ;
        RECT  0.345 1.000 0.425 1.490 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0502 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.185 0.930 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 1.635 0.600 1.965 ;
        RECT  0.085 1.220 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END CKND1

MACRO CKND12
    CLASS CORE ;
    FOREIGN CKND12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9990 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 1.060 3.095 1.450 ;
        RECT  1.850 0.345 2.935 0.655 ;
        RECT  1.350 0.345 1.850 1.450 ;
        RECT  0.685 0.345 1.350 0.655 ;
        RECT  0.325 1.060 1.350 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.6014 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 0.780 1.070 0.890 ;
        RECT  0.090 0.275 0.200 0.890 ;
        RECT  0.050 0.500 0.090 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 -0.165 3.400 0.165 ;
        RECT  3.055 -0.165 3.165 0.505 ;
        RECT  0.565 -0.165 3.055 0.165 ;
        RECT  0.455 -0.165 0.565 0.690 ;
        RECT  0.000 -0.165 0.455 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.635 3.400 1.965 ;
        RECT  0.095 1.040 0.205 1.965 ;
        RECT  0.000 1.635 0.095 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.950 1.060 3.095 1.450 ;
        RECT  1.950 0.345 2.935 0.655 ;
        RECT  0.685 0.345 1.250 0.655 ;
        RECT  0.325 1.060 1.250 1.450 ;
        RECT  2.200 0.780 3.130 0.890 ;
    END
END CKND12

MACRO CKND16
    CLASS CORE ;
    FOREIGN CKND16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.3490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.345 4.295 0.655 ;
        RECT  2.450 1.060 4.105 1.450 ;
        RECT  1.950 0.345 2.450 1.450 ;
        RECT  0.685 0.345 1.950 0.655 ;
        RECT  0.295 1.060 1.950 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.8059 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 0.780 1.670 0.890 ;
        RECT  0.090 0.275 0.200 0.890 ;
        RECT  0.050 0.500 0.090 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.565 -0.165 4.400 0.165 ;
        RECT  0.455 -0.165 0.565 0.690 ;
        RECT  0.000 -0.165 0.455 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.345 4.295 0.655 ;
        RECT  2.550 1.060 4.105 1.450 ;
        RECT  0.685 0.345 1.850 0.655 ;
        RECT  0.295 1.060 1.850 1.450 ;
        RECT  2.730 0.780 4.140 0.890 ;
    END
END CKND16

MACRO CKND2
    CLASS CORE ;
    FOREIGN CKND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.565 1.150 ;
        RECT  0.440 0.420 0.445 1.150 ;
        RECT  0.335 0.420 0.440 0.610 ;
        RECT  0.300 1.040 0.440 1.150 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1005 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.735 -0.165 0.800 0.165 ;
        RECT  0.565 -0.165 0.735 0.400 ;
        RECT  0.185 -0.165 0.565 0.165 ;
        RECT  0.075 -0.165 0.185 0.510 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 1.635 0.800 1.965 ;
        RECT  0.585 1.285 0.725 1.965 ;
        RECT  0.195 1.635 0.585 1.965 ;
        RECT  0.065 1.040 0.195 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
END CKND2

MACRO CKND20
    CLASS CORE ;
    FOREIGN CKND20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.6600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.060 5.105 1.450 ;
        RECT  2.850 0.345 4.805 0.655 ;
        RECT  2.350 0.345 2.850 1.450 ;
        RECT  0.615 0.345 2.350 0.655 ;
        RECT  0.295 1.060 2.350 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.0070 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 0.780 1.910 0.890 ;
        RECT  0.090 0.275 0.200 0.890 ;
        RECT  0.050 0.500 0.090 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.015 -0.165 5.400 0.165 ;
        RECT  4.905 -0.165 5.015 0.505 ;
        RECT  0.505 -0.165 4.905 0.165 ;
        RECT  0.395 -0.165 0.505 0.690 ;
        RECT  0.000 -0.165 0.395 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 1.060 5.105 1.450 ;
        RECT  2.950 0.345 4.805 0.655 ;
        RECT  0.615 0.345 2.250 0.655 ;
        RECT  0.295 1.060 2.250 1.450 ;
        RECT  3.260 0.780 5.140 0.890 ;
    END
END CKND20

MACRO CKND24
    CLASS CORE ;
    FOREIGN CKND24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.9920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.060 6.105 1.450 ;
        RECT  3.250 0.345 5.925 0.655 ;
        RECT  2.750 0.345 3.250 1.450 ;
        RECT  0.615 0.345 2.750 0.655 ;
        RECT  0.295 1.060 2.750 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.2090 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 0.780 2.390 0.890 ;
        RECT  0.090 0.275 0.200 0.890 ;
        RECT  0.050 0.500 0.090 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.155 -0.165 6.400 0.165 ;
        RECT  6.045 -0.165 6.155 0.505 ;
        RECT  0.505 -0.165 6.045 0.165 ;
        RECT  0.395 -0.165 0.505 0.690 ;
        RECT  0.000 -0.165 0.395 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 6.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.350 1.060 6.105 1.450 ;
        RECT  3.350 0.345 5.925 0.655 ;
        RECT  0.615 0.345 2.650 0.655 ;
        RECT  0.295 1.060 2.650 1.450 ;
        RECT  3.770 0.780 6.140 0.890 ;
    END
END CKND24

MACRO CKND2D0
    CLASS CORE ;
    FOREIGN CKND2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.290 0.755 1.150 ;
        RECT  0.555 0.290 0.645 0.400 ;
        RECT  0.455 1.040 0.645 1.150 ;
        RECT  0.345 1.040 0.455 1.470 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.555 0.930 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.165 0.800 0.165 ;
        RECT  0.085 -0.165 0.195 0.470 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.260 0.715 1.965 ;
        RECT  0.195 1.635 0.605 1.965 ;
        RECT  0.085 1.260 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END CKND2D0

MACRO CKND2D1
    CLASS CORE ;
    FOREIGN CKND2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.290 0.755 1.150 ;
        RECT  0.555 0.290 0.645 0.400 ;
        RECT  0.455 1.040 0.645 1.150 ;
        RECT  0.345 1.040 0.455 1.470 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0468 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0468 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.555 0.930 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.165 0.800 0.165 ;
        RECT  0.085 -0.165 0.195 0.580 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.260 0.715 1.965 ;
        RECT  0.195 1.635 0.605 1.965 ;
        RECT  0.085 1.040 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END CKND2D1

MACRO CKND2D2
    CLASS CORE ;
    FOREIGN CKND2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.015 1.065 1.115 ;
        RECT  0.550 0.425 0.805 0.535 ;
        RECT  0.450 0.425 0.550 1.115 ;
        RECT  0.355 1.015 0.450 1.115 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0942 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.780 1.350 1.295 ;
        RECT  1.060 0.780 1.250 0.890 ;
        RECT  0.150 1.205 1.250 1.295 ;
        RECT  0.150 0.780 0.340 0.890 ;
        RECT  0.050 0.710 0.150 1.295 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0942 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 -0.165 1.400 0.165 ;
        RECT  1.165 -0.165 1.275 0.585 ;
        RECT  0.235 -0.165 1.165 0.165 ;
        RECT  0.125 -0.165 0.235 0.585 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.400 1.965 ;
        END
    END VDD
END CKND2D2

MACRO CKND2D3
    CLASS CORE ;
    FOREIGN CKND2D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.305 1.750 1.200 ;
        RECT  0.450 0.305 1.650 0.410 ;
        RECT  1.350 1.050 1.650 1.350 ;
        RECT  0.250 1.240 1.350 1.350 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1421 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.140 ;
        RECT  0.350 1.050 1.045 1.140 ;
        RECT  0.250 0.700 0.350 1.140 ;
        RECT  0.135 0.780 0.250 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1413 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.500 1.550 0.940 ;
        RECT  0.760 0.500 1.425 0.600 ;
        RECT  0.640 0.500 0.760 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.210 -0.165 1.800 0.165 ;
        RECT  0.100 -0.165 0.210 0.555 ;
        RECT  0.000 -0.165 0.100 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.800 1.965 ;
        END
    END VDD
END CKND2D3

MACRO CKND2D4
    CLASS CORE ;
    FOREIGN CKND2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 1.050 2.250 1.350 ;
        RECT  1.890 1.050 1.950 1.270 ;
        RECT  1.800 0.475 1.890 1.270 ;
        RECT  1.585 0.475 1.800 0.585 ;
        RECT  0.540 1.180 1.800 1.270 ;
        RECT  0.540 0.475 0.755 0.585 ;
        RECT  0.450 0.475 0.540 1.270 ;
        RECT  0.445 1.105 0.450 1.270 ;
        RECT  0.335 1.105 0.445 1.525 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1874 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 0.780 2.230 0.895 ;
        RECT  1.980 0.275 2.070 0.895 ;
        RECT  1.475 0.275 1.980 0.365 ;
        RECT  1.385 0.275 1.475 0.600 ;
        RECT  1.165 0.510 1.385 0.600 ;
        RECT  1.035 0.510 1.165 0.890 ;
        RECT  0.950 0.510 1.035 0.600 ;
        RECT  0.850 0.275 0.950 0.600 ;
        RECT  0.360 0.275 0.850 0.365 ;
        RECT  0.270 0.275 0.360 0.890 ;
        RECT  0.110 0.780 0.270 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1872 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.780 1.710 0.890 ;
        RECT  1.450 0.780 1.550 1.090 ;
        RECT  0.760 0.980 1.450 1.090 ;
        RECT  0.650 0.710 0.760 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 -0.165 2.400 0.165 ;
        RECT  2.180 -0.165 2.290 0.665 ;
        RECT  1.275 -0.165 2.180 0.165 ;
        RECT  1.065 -0.165 1.275 0.415 ;
        RECT  0.180 -0.165 1.065 0.165 ;
        RECT  0.070 -0.165 0.180 0.670 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.635 2.400 1.965 ;
        RECT  2.150 1.460 2.320 1.965 ;
        RECT  1.170 1.635 2.150 1.965 ;
        RECT  1.170 1.380 1.795 1.490 ;
        RECT  1.030 1.380 1.170 1.965 ;
        RECT  0.545 1.380 1.030 1.490 ;
        RECT  0.185 1.635 1.030 1.965 ;
        RECT  0.075 1.105 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.800 0.475 1.850 1.270 ;
        RECT  1.585 0.475 1.800 0.585 ;
        RECT  0.540 1.180 1.800 1.270 ;
        RECT  0.540 0.475 0.755 0.585 ;
        RECT  0.450 0.475 0.540 1.270 ;
        RECT  0.445 1.105 0.450 1.270 ;
        RECT  0.335 1.105 0.445 1.525 ;
    END
END CKND2D4

MACRO CKND2D8
    CLASS CORE ;
    FOREIGN CKND2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.000 1.180 4.150 1.490 ;
        RECT  3.850 0.490 4.000 1.490 ;
        RECT  3.665 0.490 3.850 0.620 ;
        RECT  2.665 1.180 3.850 1.490 ;
        RECT  2.665 0.490 2.835 0.620 ;
        RECT  2.550 0.490 2.665 1.490 ;
        RECT  1.845 1.090 2.550 1.490 ;
        RECT  1.755 0.510 1.845 1.490 ;
        RECT  1.585 0.510 1.755 0.620 ;
        RECT  0.560 1.180 1.755 1.490 ;
        RECT  0.560 0.490 0.755 0.620 ;
        RECT  0.450 0.490 0.560 1.490 ;
        RECT  0.285 1.180 0.450 1.490 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.3590 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.110 0.310 4.220 0.940 ;
        RECT  3.385 0.310 4.110 0.400 ;
        RECT  3.215 0.310 3.385 0.890 ;
        RECT  2.445 0.310 3.215 0.400 ;
        RECT  2.355 0.310 2.445 0.890 ;
        RECT  2.045 0.780 2.355 0.890 ;
        RECT  1.955 0.310 2.045 0.890 ;
        RECT  1.185 0.310 1.955 0.400 ;
        RECT  1.015 0.310 1.185 0.890 ;
        RECT  0.360 0.310 1.015 0.400 ;
        RECT  0.270 0.310 0.360 0.890 ;
        RECT  0.110 0.785 0.270 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3578 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.710 1.645 0.940 ;
        RECT  1.450 0.710 1.550 1.070 ;
        RECT  0.760 0.980 1.450 1.070 ;
        RECT  0.650 0.710 0.760 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.265 -0.165 4.400 0.165 ;
        RECT  2.155 -0.165 2.265 0.620 ;
        RECT  0.180 -0.165 2.155 0.165 ;
        RECT  0.075 -0.165 0.180 0.675 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.635 4.400 1.965 ;
        RECT  0.075 1.115 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.000 1.180 4.150 1.490 ;
        RECT  3.850 0.490 4.000 1.490 ;
        RECT  3.665 0.490 3.850 0.620 ;
        RECT  2.665 1.180 3.850 1.490 ;
        RECT  2.665 0.490 2.835 0.620 ;
        RECT  2.550 0.490 2.665 1.490 ;
        RECT  1.845 1.090 1.850 1.490 ;
        RECT  1.755 0.510 1.845 1.490 ;
        RECT  1.585 0.510 1.755 0.620 ;
        RECT  0.560 1.180 1.755 1.490 ;
        RECT  0.560 0.490 0.755 0.620 ;
        RECT  0.450 0.490 0.560 1.490 ;
        RECT  0.285 1.180 0.450 1.490 ;
        RECT  3.650 0.730 3.760 1.070 ;
        RECT  2.860 0.980 3.650 1.070 ;
        RECT  2.755 0.730 2.860 1.070 ;
    END
END CKND2D8

MACRO CKND3
    CLASS CORE ;
    FOREIGN CKND3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3110 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.290 1.060 0.440 ;
        RECT  0.860 1.060 1.000 1.450 ;
        RECT  0.560 0.290 0.860 1.450 ;
        RECT  0.360 0.290 0.560 0.400 ;
        RECT  0.370 1.060 0.560 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1513 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.500 0.355 0.940 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.220 1.635 1.200 1.965 ;
        RECT  0.110 1.040 0.220 1.965 ;
        RECT  0.000 1.635 0.110 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.290 1.060 0.440 ;
        RECT  0.950 1.060 1.000 1.450 ;
        RECT  0.360 0.290 0.450 0.400 ;
        RECT  0.370 1.060 0.450 1.450 ;
    END
END CKND3

MACRO CKND4
    CLASS CORE ;
    FOREIGN CKND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.335 1.075 0.595 ;
        RECT  0.850 1.060 1.075 1.450 ;
        RECT  0.550 0.335 0.850 1.450 ;
        RECT  0.385 0.335 0.550 0.595 ;
        RECT  0.385 1.060 0.550 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2010 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 -0.165 1.400 0.165 ;
        RECT  1.195 -0.165 1.305 0.545 ;
        RECT  0.265 -0.165 1.195 0.165 ;
        RECT  0.155 -0.165 0.265 0.545 ;
        RECT  0.000 -0.165 0.155 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 1.635 1.400 1.965 ;
        RECT  1.195 1.040 1.305 1.965 ;
        RECT  0.265 1.635 1.195 1.965 ;
        RECT  0.155 1.260 0.265 1.965 ;
        RECT  0.000 1.635 0.155 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.335 1.075 0.595 ;
        RECT  0.950 1.060 1.075 1.450 ;
        RECT  0.385 0.335 0.450 0.595 ;
        RECT  0.385 1.060 0.450 1.450 ;
    END
END CKND4

MACRO CKND6
    CLASS CORE ;
    FOREIGN CKND6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.345 1.525 0.655 ;
        RECT  1.250 1.060 1.505 1.450 ;
        RECT  0.950 0.345 1.250 1.450 ;
        RECT  0.335 0.345 0.950 0.655 ;
        RECT  0.295 1.060 0.950 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.3017 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 0.780 0.750 0.890 ;
        RECT  0.090 0.275 0.200 0.890 ;
        RECT  0.050 0.500 0.090 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.345 1.525 0.655 ;
        RECT  1.350 1.060 1.505 1.450 ;
        RECT  0.335 0.345 0.850 0.655 ;
        RECT  0.295 1.060 0.850 1.450 ;
    END
END CKND6

MACRO CKND8
    CLASS CORE ;
    FOREIGN CKND8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6810 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.345 2.355 0.655 ;
        RECT  1.450 1.060 2.055 1.450 ;
        RECT  0.950 0.345 1.450 1.450 ;
        RECT  0.685 0.345 0.950 0.655 ;
        RECT  0.325 1.060 0.950 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.4011 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 0.780 0.670 0.890 ;
        RECT  0.090 0.275 0.200 0.890 ;
        RECT  0.050 0.500 0.090 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.565 -0.165 2.400 0.165 ;
        RECT  0.455 -0.165 0.565 0.690 ;
        RECT  0.000 -0.165 0.455 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.285 1.635 2.400 1.965 ;
        RECT  2.175 1.040 2.285 1.965 ;
        RECT  0.205 1.635 2.175 1.965 ;
        RECT  0.095 1.040 0.205 1.965 ;
        RECT  0.000 1.635 0.095 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.550 0.345 2.355 0.655 ;
        RECT  1.550 1.060 2.055 1.450 ;
        RECT  0.685 0.345 0.850 0.655 ;
        RECT  0.325 1.060 0.850 1.450 ;
        RECT  1.720 0.780 2.130 0.890 ;
    END
END CKND8

MACRO CKXOR2D0
    CLASS CORE ;
    FOREIGN CKXOR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.310 1.950 1.490 ;
        RECT  1.820 0.310 1.850 0.695 ;
        RECT  1.820 1.240 1.850 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0259 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.405 0.700 1.450 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0510 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.165 2.000 0.165 ;
        RECT  0.320 -0.165 0.510 0.385 ;
        RECT  0.000 -0.165 0.320 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.475 1.635 2.000 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.730 0.770 1.760 0.940 ;
        RECT  1.640 0.305 1.730 1.495 ;
        RECT  0.880 0.305 1.640 0.405 ;
        RECT  0.935 1.390 1.640 1.495 ;
        RECT  1.315 1.210 1.430 1.300 ;
        RECT  1.215 0.495 1.315 1.300 ;
        RECT  0.705 1.210 1.215 1.300 ;
        RECT  1.015 0.545 1.105 1.120 ;
        RECT  0.595 0.545 1.015 0.655 ;
        RECT  0.650 1.020 1.015 1.120 ;
        RECT  0.370 0.790 0.925 0.900 ;
        RECT  0.595 1.210 0.705 1.525 ;
        RECT  0.280 0.510 0.370 1.290 ;
        RECT  0.185 0.510 0.280 0.600 ;
        RECT  0.185 1.200 0.280 1.290 ;
        RECT  0.075 0.370 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.490 ;
    END
END CKXOR2D0

MACRO CKXOR2D1
    CLASS CORE ;
    FOREIGN CKXOR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.275 1.950 1.490 ;
        RECT  1.820 0.275 1.850 0.675 ;
        RECT  1.820 1.045 1.850 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.405 0.700 1.450 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0582 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.165 2.000 0.165 ;
        RECT  0.320 -0.165 0.510 0.385 ;
        RECT  0.000 -0.165 0.320 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.475 1.635 2.000 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.730 0.750 1.760 0.920 ;
        RECT  1.640 0.305 1.730 1.495 ;
        RECT  0.880 0.305 1.640 0.405 ;
        RECT  0.935 1.390 1.640 1.495 ;
        RECT  1.315 1.210 1.430 1.300 ;
        RECT  1.215 0.495 1.315 1.300 ;
        RECT  0.705 1.210 1.215 1.300 ;
        RECT  1.015 0.520 1.105 1.120 ;
        RECT  0.595 0.520 1.015 0.630 ;
        RECT  0.650 1.020 1.015 1.120 ;
        RECT  0.370 0.790 0.925 0.900 ;
        RECT  0.595 1.210 0.705 1.525 ;
        RECT  0.280 0.510 0.370 1.290 ;
        RECT  0.185 0.510 0.280 0.600 ;
        RECT  0.185 1.200 0.280 1.290 ;
        RECT  0.075 0.390 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.490 ;
    END
END CKXOR2D1

MACRO CKXOR2D2
    CLASS CORE ;
    FOREIGN CKXOR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.310 1.950 1.505 ;
        RECT  1.700 0.310 1.850 0.420 ;
        RECT  1.725 1.395 1.850 1.505 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.405 0.700 1.450 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0735 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.165 2.200 0.165 ;
        RECT  0.320 -0.165 0.510 0.385 ;
        RECT  0.000 -0.165 0.320 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.475 1.635 2.200 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.660 0.510 1.760 1.290 ;
        RECT  1.590 0.510 1.660 0.610 ;
        RECT  1.635 1.190 1.660 1.290 ;
        RECT  1.535 1.190 1.635 1.495 ;
        RECT  1.490 0.305 1.590 0.610 ;
        RECT  0.930 1.390 1.535 1.495 ;
        RECT  0.880 0.305 1.490 0.405 ;
        RECT  1.315 1.210 1.425 1.300 ;
        RECT  1.215 0.495 1.315 1.300 ;
        RECT  0.700 1.210 1.215 1.300 ;
        RECT  1.015 0.520 1.105 1.120 ;
        RECT  0.595 0.520 1.015 0.630 ;
        RECT  0.645 1.020 1.015 1.120 ;
        RECT  0.370 0.790 0.920 0.900 ;
        RECT  0.590 1.210 0.700 1.525 ;
        RECT  0.280 0.510 0.370 1.290 ;
        RECT  0.185 0.510 0.280 0.600 ;
        RECT  0.185 1.200 0.280 1.290 ;
        RECT  0.075 0.390 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.460 ;
    END
END CKXOR2D2

MACRO CKXOR2D4
    CLASS CORE ;
    FOREIGN CKXOR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.755 0.275 3.865 0.705 ;
        RECT  3.755 1.030 3.865 1.480 ;
        RECT  3.650 0.595 3.755 0.705 ;
        RECT  3.650 1.030 3.755 1.140 ;
        RECT  3.365 0.595 3.650 1.140 ;
        RECT  3.350 0.595 3.365 1.490 ;
        RECT  3.345 0.595 3.350 0.705 ;
        RECT  3.250 1.030 3.350 1.490 ;
        RECT  3.235 0.275 3.345 0.705 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.355 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1418 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.700 2.950 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.665 ;
        RECT  3.605 -0.165 4.015 0.165 ;
        RECT  3.495 -0.165 3.605 0.495 ;
        RECT  0.000 -0.165 3.495 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.135 4.125 1.965 ;
        RECT  3.110 1.635 4.015 1.965 ;
        RECT  2.940 1.455 3.110 1.965 ;
        RECT  0.000 1.635 2.940 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.755 0.275 3.865 0.705 ;
        RECT  3.755 1.030 3.865 1.480 ;
        RECT  3.750 0.595 3.755 0.705 ;
        RECT  3.750 1.030 3.755 1.140 ;
        RECT  3.235 0.275 3.250 0.705 ;
        RECT  3.040 0.325 3.145 1.345 ;
        RECT  2.470 0.325 3.040 0.425 ;
        RECT  2.535 1.255 3.040 1.345 ;
        RECT  2.550 1.035 2.845 1.145 ;
        RECT  2.550 0.515 2.820 0.610 ;
        RECT  2.440 0.515 2.550 1.145 ;
        RECT  2.425 1.255 2.535 1.495 ;
        RECT  2.370 0.275 2.470 0.425 ;
        RECT  1.990 0.275 2.370 0.365 ;
        RECT  2.280 0.655 2.335 1.185 ;
        RECT  2.275 0.455 2.280 1.185 ;
        RECT  2.245 0.455 2.275 1.525 ;
        RECT  2.110 0.455 2.245 0.750 ;
        RECT  2.165 1.085 2.245 1.525 ;
        RECT  0.685 1.435 2.165 1.525 ;
        RECT  1.955 0.875 2.155 0.975 ;
        RECT  1.905 1.065 2.015 1.345 ;
        RECT  1.880 0.275 1.990 0.545 ;
        RECT  1.845 0.660 1.955 0.975 ;
        RECT  1.380 1.065 1.905 1.160 ;
        RECT  1.380 0.455 1.880 0.545 ;
        RECT  1.490 0.660 1.845 0.760 ;
        RECT  1.200 1.255 1.795 1.345 ;
        RECT  1.200 0.275 1.770 0.365 ;
        RECT  1.290 0.455 1.380 1.160 ;
        RECT  1.110 0.275 1.200 1.345 ;
        RECT  1.075 0.275 1.110 0.590 ;
        RECT  1.075 1.090 1.110 1.345 ;
        RECT  0.685 0.750 1.020 0.920 ;
        RECT  0.575 0.275 0.685 1.525 ;
        RECT  0.185 0.510 0.575 0.600 ;
        RECT  0.185 1.435 0.575 1.525 ;
        RECT  0.075 0.360 0.185 0.600 ;
        RECT  0.075 1.210 0.185 1.525 ;
    END
END CKXOR2D4

MACRO CMPE42D1
    CLASS CORE ;
    FOREIGN CMPE42D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.050 0.275 9.150 1.490 ;
        RECT  9.015 0.275 9.050 0.665 ;
        RECT  9.020 1.040 9.050 1.490 ;
        END
    END S
    PIN D
        ANTENNAGATEAREA 0.0952 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.510 6.350 0.920 ;
        RECT  6.110 0.750 6.250 0.920 ;
        END
    END D
    PIN COX
        ANTENNADIFFAREA 0.1420 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.750 0.325 4.785 0.645 ;
        RECT  4.665 0.325 4.750 1.165 ;
        RECT  4.645 0.510 4.665 1.165 ;
        RECT  4.605 0.995 4.645 1.165 ;
        END
    END COX
    PIN CO
        ANTENNADIFFAREA 0.1400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.645 0.310 8.750 0.690 ;
        RECT  8.630 0.510 8.645 0.690 ;
        RECT  8.450 0.510 8.630 1.150 ;
        END
    END CO
    PIN CIX
        ANTENNAGATEAREA 0.0529 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.230 0.510 8.350 0.890 ;
        RECT  8.165 0.710 8.230 0.890 ;
        END
    END CIX
    PIN C
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.425 0.510 4.555 0.890 ;
        RECT  4.340 0.710 4.425 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0669 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.195 0.700 1.350 1.100 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.440 0.895 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 9.200 0.165 ;
        RECT  0.075 -0.165 0.185 0.475 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.635 9.200 1.965 ;
        RECT  0.075 1.325 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.880 0.775 8.960 0.945 ;
        RECT  8.780 0.775 8.880 1.345 ;
        RECT  7.570 1.255 8.780 1.345 ;
        RECT  7.285 1.435 8.525 1.525 ;
        RECT  8.075 0.275 8.455 0.410 ;
        RECT  8.075 0.980 8.360 1.150 ;
        RECT  7.985 0.275 8.075 1.150 ;
        RECT  7.375 0.275 7.985 0.365 ;
        RECT  7.905 0.720 7.985 0.890 ;
        RECT  7.815 0.455 7.895 0.625 ;
        RECT  7.815 0.995 7.845 1.165 ;
        RECT  7.725 0.455 7.815 1.165 ;
        RECT  7.675 0.995 7.725 1.165 ;
        RECT  7.570 0.465 7.635 0.635 ;
        RECT  7.475 0.465 7.570 1.345 ;
        RECT  7.400 1.145 7.475 1.345 ;
        RECT  7.285 0.275 7.375 0.975 ;
        RECT  7.250 0.275 7.285 1.300 ;
        RECT  7.065 1.420 7.285 1.525 ;
        RECT  7.175 0.885 7.250 1.300 ;
        RECT  7.065 0.440 7.140 0.635 ;
        RECT  6.965 0.440 7.065 1.525 ;
        RECT  6.885 1.420 6.965 1.525 ;
        RECT  6.770 0.475 6.875 1.330 ;
        RECT  5.545 0.275 6.785 0.365 ;
        RECT  6.760 0.475 6.770 1.525 ;
        RECT  6.640 1.240 6.760 1.525 ;
        RECT  6.555 0.530 6.670 1.145 ;
        RECT  6.015 1.240 6.640 1.335 ;
        RECT  6.445 0.530 6.555 0.670 ;
        RECT  6.385 1.035 6.555 1.145 ;
        RECT  6.015 0.555 6.140 0.655 ;
        RECT  5.925 0.555 6.015 1.505 ;
        RECT  5.885 0.775 5.925 1.505 ;
        RECT  5.830 0.775 5.885 0.945 ;
        RECT  5.740 0.455 5.830 0.625 ;
        RECT  5.740 1.060 5.755 1.525 ;
        RECT  5.635 0.455 5.740 1.525 ;
        RECT  4.975 1.435 5.635 1.525 ;
        RECT  5.440 0.275 5.545 1.330 ;
        RECT  5.405 1.160 5.440 1.330 ;
        RECT  5.235 0.325 5.310 1.065 ;
        RECT  5.220 0.325 5.235 1.330 ;
        RECT  5.195 0.325 5.220 0.580 ;
        RECT  5.125 0.975 5.220 1.330 ;
        RECT  4.975 0.715 5.130 0.885 ;
        RECT  4.885 0.715 4.975 1.525 ;
        RECT  3.695 1.255 4.885 1.345 ;
        RECT  3.205 1.435 4.665 1.525 ;
        RECT  4.215 0.275 4.575 0.420 ;
        RECT  4.215 1.000 4.515 1.155 ;
        RECT  4.125 0.275 4.215 1.155 ;
        RECT  3.515 0.275 4.125 0.365 ;
        RECT  4.045 0.735 4.125 0.905 ;
        RECT  3.955 0.465 4.035 0.635 ;
        RECT  3.955 1.020 3.995 1.165 ;
        RECT  3.865 0.465 3.955 1.165 ;
        RECT  3.805 1.020 3.865 1.165 ;
        RECT  3.695 0.455 3.775 0.640 ;
        RECT  3.605 0.455 3.695 1.345 ;
        RECT  3.555 1.105 3.605 1.345 ;
        RECT  3.430 0.275 3.515 0.920 ;
        RECT  3.415 0.275 3.430 1.275 ;
        RECT  3.325 0.790 3.415 1.275 ;
        RECT  3.055 0.425 3.205 1.525 ;
        RECT  2.865 0.470 2.955 1.450 ;
        RECT  2.840 0.470 2.865 0.640 ;
        RECT  2.170 1.320 2.865 1.450 ;
        RECT  2.720 0.745 2.775 0.915 ;
        RECT  2.630 0.360 2.720 1.185 ;
        RECT  2.600 0.360 2.630 0.595 ;
        RECT  2.495 1.075 2.630 1.185 ;
        RECT  2.480 0.750 2.540 0.920 ;
        RECT  2.390 0.275 2.480 0.920 ;
        RECT  1.665 0.275 2.390 0.365 ;
        RECT  2.170 0.475 2.260 0.675 ;
        RECT  2.060 0.475 2.170 1.450 ;
        RECT  2.035 0.775 2.060 1.450 ;
        RECT  1.970 0.775 2.035 0.945 ;
        RECT  1.865 0.465 1.950 0.655 ;
        RECT  1.865 1.070 1.925 1.525 ;
        RECT  1.775 0.465 1.865 1.525 ;
        RECT  0.680 1.435 1.775 1.525 ;
        RECT  1.555 0.275 1.665 1.325 ;
        RECT  1.090 1.210 1.445 1.320 ;
        RECT  1.295 0.340 1.405 0.610 ;
        RECT  1.090 0.500 1.295 0.610 ;
        RECT  1.000 0.500 1.090 1.320 ;
        RECT  0.945 0.500 1.000 0.675 ;
        RECT  0.790 1.210 1.000 1.320 ;
        RECT  0.830 0.275 0.945 0.675 ;
        RECT  0.680 0.780 0.890 0.895 ;
        RECT  0.590 0.575 0.680 1.525 ;
        RECT  0.445 0.575 0.590 0.675 ;
        RECT  0.445 1.435 0.590 1.525 ;
        RECT  0.335 0.275 0.445 0.675 ;
        RECT  0.335 1.025 0.445 1.525 ;
    END
END CMPE42D1

MACRO CMPE42D2
    CLASS CORE ;
    FOREIGN CMPE42D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.050 0.275 9.175 1.295 ;
        END
    END S
    PIN D
        ANTENNAGATEAREA 0.0945 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.700 6.550 1.100 ;
        RECT  6.280 0.790 6.450 0.890 ;
        END
    END D
    PIN COX
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.950 1.000 4.985 1.095 ;
        RECT  4.850 0.310 4.950 1.095 ;
        RECT  4.805 0.310 4.850 0.600 ;
        RECT  4.795 1.000 4.850 1.095 ;
        END
    END COX
    PIN CO
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.650 0.275 9.750 1.490 ;
        RECT  9.565 0.275 9.650 0.685 ;
        RECT  9.570 1.040 9.650 1.490 ;
        END
    END CO
    PIN CIX
        ANTENNAGATEAREA 0.0529 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.645 0.510 8.755 0.900 ;
        RECT  8.550 0.780 8.645 0.900 ;
        END
    END CIX
    PIN C
        ANTENNAGATEAREA 0.0529 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.710 4.750 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.350 1.100 ;
        RECT  1.195 0.700 1.250 0.920 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.440 0.895 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.555 -0.165 10.000 0.165 ;
        RECT  6.385 -0.165 6.555 0.285 ;
        RECT  5.175 -0.165 6.385 0.165 ;
        RECT  5.065 -0.165 5.175 0.550 ;
        RECT  0.185 -0.165 5.065 0.165 ;
        RECT  0.075 -0.165 0.185 0.475 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.540 1.635 10.000 1.965 ;
        RECT  6.370 1.445 6.540 1.965 ;
        RECT  0.185 1.635 6.370 1.965 ;
        RECT  0.075 1.325 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.450 0.780 9.560 0.890 ;
        RECT  9.350 0.780 9.450 1.475 ;
        RECT  7.285 1.385 9.350 1.475 ;
        RECT  8.935 0.730 8.960 0.940 ;
        RECT  8.845 0.730 8.935 1.295 ;
        RECT  7.850 1.205 8.845 1.295 ;
        RECT  8.420 0.275 8.745 0.420 ;
        RECT  8.420 1.015 8.735 1.115 ;
        RECT  8.330 0.275 8.420 1.115 ;
        RECT  7.660 0.275 8.330 0.365 ;
        RECT  8.220 0.750 8.330 0.920 ;
        RECT  8.130 0.495 8.240 0.605 ;
        RECT  8.040 0.495 8.130 1.115 ;
        RECT  7.960 1.015 8.040 1.115 ;
        RECT  7.850 0.455 7.930 0.865 ;
        RECT  7.820 0.455 7.850 1.295 ;
        RECT  7.760 0.775 7.820 1.295 ;
        RECT  7.655 1.185 7.760 1.295 ;
        RECT  7.550 0.275 7.660 1.055 ;
        RECT  7.545 0.965 7.550 1.055 ;
        RECT  7.435 0.965 7.545 1.255 ;
        RECT  7.290 0.440 7.400 0.875 ;
        RECT  7.285 0.775 7.290 0.875 ;
        RECT  7.175 0.775 7.285 1.475 ;
        RECT  7.065 0.525 7.165 0.635 ;
        RECT  7.025 0.525 7.065 1.340 ;
        RECT  6.825 0.275 7.060 0.375 ;
        RECT  6.975 0.525 7.025 1.525 ;
        RECT  6.915 1.250 6.975 1.525 ;
        RECT  6.215 1.250 6.915 1.340 ;
        RECT  6.785 0.555 6.885 1.140 ;
        RECT  6.735 0.275 6.825 0.465 ;
        RECT  6.650 0.555 6.785 0.655 ;
        RECT  6.660 1.030 6.785 1.140 ;
        RECT  6.275 0.375 6.735 0.465 ;
        RECT  6.190 0.555 6.290 0.655 ;
        RECT  6.185 0.275 6.275 0.465 ;
        RECT  6.190 1.035 6.215 1.495 ;
        RECT  6.100 0.555 6.190 1.495 ;
        RECT  5.695 0.275 6.185 0.365 ;
        RECT  6.025 0.775 6.100 0.945 ;
        RECT  5.915 0.535 6.010 0.645 ;
        RECT  5.915 1.060 5.960 1.525 ;
        RECT  5.825 0.535 5.915 1.525 ;
        RECT  5.190 1.435 5.825 1.525 ;
        RECT  5.585 0.275 5.695 1.330 ;
        RECT  5.375 0.340 5.465 1.330 ;
        RECT  5.330 0.340 5.375 0.550 ;
        RECT  5.325 1.120 5.375 1.330 ;
        RECT  5.190 0.715 5.270 0.885 ;
        RECT  5.100 0.715 5.190 1.525 ;
        RECT  3.800 1.185 5.100 1.275 ;
        RECT  4.630 1.365 4.840 1.525 ;
        RECT  4.320 0.275 4.695 0.420 ;
        RECT  4.320 1.000 4.685 1.095 ;
        RECT  3.235 1.365 4.630 1.455 ;
        RECT  4.230 0.275 4.320 1.095 ;
        RECT  3.610 0.275 4.230 0.365 ;
        RECT  4.170 0.735 4.230 0.905 ;
        RECT  4.080 0.455 4.140 0.625 ;
        RECT  3.990 0.455 4.080 1.095 ;
        RECT  3.910 0.985 3.990 1.095 ;
        RECT  3.800 0.455 3.880 0.640 ;
        RECT  3.710 0.455 3.800 1.275 ;
        RECT  3.605 1.165 3.710 1.275 ;
        RECT  3.500 0.275 3.610 0.920 ;
        RECT  3.495 0.790 3.500 0.920 ;
        RECT  3.385 0.790 3.495 1.275 ;
        RECT  3.235 0.490 3.390 0.600 ;
        RECT  3.125 0.490 3.235 1.455 ;
        RECT  2.975 0.475 3.035 1.340 ;
        RECT  2.940 0.475 2.975 1.465 ;
        RECT  2.865 1.250 2.940 1.465 ;
        RECT  2.200 1.250 2.865 1.340 ;
        RECT  2.745 0.575 2.850 1.135 ;
        RECT  2.740 0.275 2.745 1.135 ;
        RECT  2.635 0.275 2.740 0.675 ;
        RECT  2.550 1.025 2.740 1.135 ;
        RECT  2.495 0.780 2.615 0.890 ;
        RECT  2.405 0.275 2.495 0.890 ;
        RECT  1.680 0.275 2.405 0.365 ;
        RECT  2.200 0.545 2.255 0.645 ;
        RECT  2.085 0.545 2.200 1.340 ;
        RECT  2.010 0.775 2.085 0.945 ;
        RECT  1.900 0.465 1.955 0.655 ;
        RECT  1.900 1.045 1.945 1.525 ;
        RECT  1.810 0.465 1.900 1.525 ;
        RECT  0.680 1.435 1.810 1.525 ;
        RECT  1.570 0.275 1.680 1.325 ;
        RECT  1.090 1.210 1.460 1.320 ;
        RECT  1.310 0.340 1.420 0.590 ;
        RECT  1.090 0.500 1.310 0.590 ;
        RECT  1.000 0.500 1.090 1.320 ;
        RECT  0.945 0.500 1.000 0.675 ;
        RECT  0.790 1.210 1.000 1.320 ;
        RECT  0.830 0.275 0.945 0.675 ;
        RECT  0.680 0.780 0.890 0.895 ;
        RECT  0.590 0.575 0.680 1.525 ;
        RECT  0.445 0.575 0.590 0.675 ;
        RECT  0.445 1.435 0.590 1.525 ;
        RECT  0.335 0.275 0.445 0.675 ;
        RECT  0.335 1.025 0.445 1.525 ;
    END
END CMPE42D2

MACRO DCAP
    CLASS CORE ;
    FOREIGN DCAP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.215 -0.165 0.600 0.165 ;
        RECT  0.105 -0.165 0.215 0.530 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.635 0.600 1.965 ;
        RECT  0.115 1.330 0.225 1.965 ;
        RECT  0.000 1.635 0.115 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.475 0.810 0.530 1.020 ;
        RECT  0.375 1.110 0.485 1.540 ;
        RECT  0.365 0.335 0.475 1.020 ;
        RECT  0.200 1.110 0.375 1.220 ;
        RECT  0.090 0.620 0.200 1.220 ;
    END
END DCAP

MACRO DCAP16
    CLASS CORE ;
    FOREIGN DCAP16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.865 -0.165 3.200 0.165 ;
        RECT  2.755 -0.165 2.865 0.555 ;
        RECT  1.965 -0.165 2.755 0.165 ;
        RECT  1.855 -0.165 1.965 0.555 ;
        RECT  1.075 -0.165 1.855 0.165 ;
        RECT  0.965 -0.165 1.075 0.555 ;
        RECT  0.185 -0.165 0.965 0.165 ;
        RECT  0.075 -0.165 0.185 0.555 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.865 1.635 3.200 1.965 ;
        RECT  2.755 1.335 2.865 1.965 ;
        RECT  1.965 1.635 2.755 1.965 ;
        RECT  1.855 1.085 1.965 1.965 ;
        RECT  1.075 1.635 1.855 1.965 ;
        RECT  0.965 1.085 1.075 1.965 ;
        RECT  0.185 1.635 0.965 1.965 ;
        RECT  0.075 1.070 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.015 0.345 3.125 1.065 ;
        RECT  3.015 1.155 3.125 1.390 ;
        RECT  2.910 0.950 3.015 1.065 ;
        RECT  2.800 1.155 3.015 1.245 ;
        RECT  2.690 0.645 2.800 1.245 ;
        RECT  0.385 0.645 2.690 0.755 ;
    END
END DCAP16

MACRO DCAP32
    CLASS CORE ;
    FOREIGN DCAP32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.065 -0.165 6.400 0.165 ;
        RECT  5.955 -0.165 6.065 0.555 ;
        RECT  4.885 -0.165 5.955 0.165 ;
        RECT  4.775 -0.165 4.885 0.555 ;
        RECT  3.710 -0.165 4.775 0.165 ;
        RECT  3.600 -0.165 3.710 0.555 ;
        RECT  2.535 -0.165 3.600 0.165 ;
        RECT  2.425 -0.165 2.535 0.555 ;
        RECT  1.360 -0.165 2.425 0.165 ;
        RECT  1.250 -0.165 1.360 0.555 ;
        RECT  0.185 -0.165 1.250 0.165 ;
        RECT  0.075 -0.165 0.185 0.555 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.065 1.635 6.400 1.965 ;
        RECT  5.955 1.335 6.065 1.965 ;
        RECT  4.895 1.635 5.955 1.965 ;
        RECT  4.765 1.085 4.895 1.965 ;
        RECT  3.720 1.635 4.765 1.965 ;
        RECT  3.590 1.085 3.720 1.965 ;
        RECT  2.545 1.635 3.590 1.965 ;
        RECT  2.415 1.085 2.545 1.965 ;
        RECT  1.370 1.635 2.415 1.965 ;
        RECT  1.240 1.085 1.370 1.965 ;
        RECT  0.195 1.635 1.240 1.965 ;
        RECT  0.065 1.085 0.195 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.215 0.345 6.325 1.065 ;
        RECT  6.215 1.155 6.325 1.390 ;
        RECT  6.110 0.950 6.215 1.065 ;
        RECT  5.910 1.155 6.215 1.245 ;
        RECT  5.800 0.645 5.910 1.245 ;
        RECT  0.385 0.645 5.800 0.755 ;
    END
END DCAP32

MACRO DCAP4
    CLASS CORE ;
    FOREIGN DCAP4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.465 -0.165 0.800 0.165 ;
        RECT  0.355 -0.165 0.465 0.555 ;
        RECT  0.185 -0.165 0.355 0.165 ;
        RECT  0.075 -0.165 0.185 0.555 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.465 1.635 0.800 1.965 ;
        RECT  0.355 1.325 0.465 1.965 ;
        RECT  0.185 1.635 0.355 1.965 ;
        RECT  0.075 1.070 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.615 0.345 0.725 0.995 ;
        RECT  0.615 1.105 0.725 1.390 ;
        RECT  0.510 0.880 0.615 0.995 ;
        RECT  0.405 1.105 0.615 1.215 ;
        RECT  0.295 0.675 0.405 1.215 ;
        RECT  0.100 0.675 0.295 0.785 ;
    END
END DCAP4

MACRO DCAP64
    CLASS CORE ;
    FOREIGN DCAP64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.465 -0.165 12.800 0.165 ;
        RECT  12.355 -0.165 12.465 0.555 ;
        RECT  11.335 -0.165 12.355 0.165 ;
        RECT  11.225 -0.165 11.335 0.555 ;
        RECT  10.220 -0.165 11.225 0.165 ;
        RECT  10.110 -0.165 10.220 0.555 ;
        RECT  9.105 -0.165 10.110 0.165 ;
        RECT  8.995 -0.165 9.105 0.555 ;
        RECT  7.990 -0.165 8.995 0.165 ;
        RECT  7.880 -0.165 7.990 0.555 ;
        RECT  6.875 -0.165 7.880 0.165 ;
        RECT  6.765 -0.165 6.875 0.555 ;
        RECT  5.760 -0.165 6.765 0.165 ;
        RECT  5.650 -0.165 5.760 0.555 ;
        RECT  4.645 -0.165 5.650 0.165 ;
        RECT  4.535 -0.165 4.645 0.555 ;
        RECT  3.530 -0.165 4.535 0.165 ;
        RECT  3.420 -0.165 3.530 0.555 ;
        RECT  2.415 -0.165 3.420 0.165 ;
        RECT  2.305 -0.165 2.415 0.555 ;
        RECT  1.300 -0.165 2.305 0.165 ;
        RECT  1.190 -0.165 1.300 0.555 ;
        RECT  0.185 -0.165 1.190 0.165 ;
        RECT  0.075 -0.165 0.185 0.555 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.465 1.635 12.800 1.965 ;
        RECT  12.355 1.335 12.465 1.965 ;
        RECT  11.345 1.635 12.355 1.965 ;
        RECT  11.215 1.085 11.345 1.965 ;
        RECT  10.230 1.635 11.215 1.965 ;
        RECT  10.100 1.085 10.230 1.965 ;
        RECT  9.115 1.635 10.100 1.965 ;
        RECT  8.985 1.085 9.115 1.965 ;
        RECT  8.000 1.635 8.985 1.965 ;
        RECT  7.870 1.085 8.000 1.965 ;
        RECT  6.885 1.635 7.870 1.965 ;
        RECT  6.755 1.085 6.885 1.965 ;
        RECT  5.770 1.635 6.755 1.965 ;
        RECT  5.640 1.085 5.770 1.965 ;
        RECT  4.655 1.635 5.640 1.965 ;
        RECT  4.525 1.085 4.655 1.965 ;
        RECT  3.540 1.635 4.525 1.965 ;
        RECT  3.410 1.085 3.540 1.965 ;
        RECT  2.425 1.635 3.410 1.965 ;
        RECT  2.295 1.085 2.425 1.965 ;
        RECT  1.310 1.635 2.295 1.965 ;
        RECT  1.180 1.085 1.310 1.965 ;
        RECT  0.185 1.635 1.180 1.965 ;
        RECT  0.075 1.070 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  12.615 0.345 12.725 1.065 ;
        RECT  12.615 1.155 12.725 1.390 ;
        RECT  12.510 0.950 12.615 1.065 ;
        RECT  12.310 1.155 12.615 1.245 ;
        RECT  12.200 0.645 12.310 1.245 ;
        RECT  0.305 0.645 12.200 0.755 ;
    END
END DCAP64

MACRO DCAP8
    CLASS CORE ;
    FOREIGN DCAP8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 -0.165 1.600 0.165 ;
        RECT  1.155 -0.165 1.265 0.555 ;
        RECT  0.185 -0.165 1.155 0.165 ;
        RECT  0.075 -0.165 0.185 0.555 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 1.635 1.600 1.965 ;
        RECT  1.155 1.335 1.265 1.965 ;
        RECT  0.185 1.635 1.155 1.965 ;
        RECT  0.075 1.070 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.415 0.345 1.525 1.065 ;
        RECT  1.415 1.155 1.525 1.390 ;
        RECT  1.310 0.950 1.415 1.065 ;
        RECT  1.200 1.155 1.415 1.245 ;
        RECT  1.090 0.645 1.200 1.245 ;
        RECT  0.240 0.645 1.090 0.755 ;
    END
END DCAP8

MACRO DEL0
    CLASS CORE ;
    FOREIGN DEL0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.280 2.550 1.490 ;
        RECT  2.415 0.280 2.450 0.490 ;
        RECT  2.415 1.280 2.450 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.940 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 0.585 2.360 1.150 ;
        RECT  1.485 0.585 2.260 0.695 ;
        RECT  1.485 1.040 2.260 1.150 ;
        RECT  1.225 0.785 1.985 0.890 ;
        RECT  1.375 0.275 1.485 0.695 ;
        RECT  1.375 1.040 1.485 1.470 ;
        RECT  1.115 0.275 1.225 1.470 ;
        RECT  0.585 0.780 0.905 0.890 ;
        RECT  0.475 0.500 0.585 1.150 ;
        RECT  0.185 0.500 0.475 0.600 ;
        RECT  0.185 1.050 0.475 1.150 ;
        RECT  0.075 0.350 0.185 0.600 ;
        RECT  0.075 1.050 0.185 1.480 ;
    END
END DEL0

MACRO DEL005
    CLASS CORE ;
    FOREIGN DEL005 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.065 0.510 1.150 1.090 ;
        RECT  1.050 0.510 1.065 1.485 ;
        RECT  0.935 0.275 1.050 0.675 ;
        RECT  0.935 0.990 1.050 1.485 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.755 0.555 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.780 -0.165 1.200 0.165 ;
        RECT  0.610 -0.165 0.780 0.285 ;
        RECT  0.000 -0.165 0.610 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.765 1.635 1.200 1.965 ;
        RECT  0.645 1.040 0.765 1.965 ;
        RECT  0.000 1.635 0.645 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.715 0.375 0.825 0.940 ;
        RECT  0.185 0.375 0.715 0.465 ;
        RECT  0.355 0.555 0.515 0.655 ;
        RECT  0.355 1.380 0.515 1.490 ;
        RECT  0.265 0.555 0.355 1.490 ;
        RECT  0.175 0.275 0.185 0.465 ;
        RECT  0.075 0.275 0.175 1.470 ;
    END
END DEL005

MACRO DEL01
    CLASS CORE ;
    FOREIGN DEL01 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.310 2.150 1.490 ;
        RECT  1.970 0.310 2.050 0.520 ;
        RECT  2.015 1.040 2.050 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.200 0.710 0.250 0.940 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.860 -0.165 2.200 0.165 ;
        RECT  1.705 -0.165 1.860 0.620 ;
        RECT  0.505 -0.165 1.705 0.165 ;
        RECT  0.335 -0.165 0.505 0.410 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.635 2.200 1.965 ;
        RECT  1.700 1.465 1.870 1.965 ;
        RECT  0.505 1.635 1.700 1.965 ;
        RECT  0.335 1.390 0.505 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.855 0.730 1.960 0.940 ;
        RECT  1.725 0.730 1.855 1.375 ;
        RECT  1.335 1.285 1.725 1.375 ;
        RECT  1.445 0.275 1.555 1.195 ;
        RECT  1.295 0.540 1.335 1.375 ;
        RECT  1.245 0.275 1.295 1.470 ;
        RECT  1.185 0.275 1.245 0.695 ;
        RECT  1.185 1.030 1.245 1.470 ;
        RECT  1.000 0.785 1.155 0.895 ;
        RECT  0.890 0.275 1.000 1.470 ;
        RECT  0.740 0.540 0.800 1.140 ;
        RECT  0.710 0.275 0.740 1.470 ;
        RECT  0.630 0.275 0.710 0.695 ;
        RECT  0.630 1.040 0.710 1.470 ;
        RECT  0.540 0.785 0.620 0.895 ;
        RECT  0.450 0.500 0.540 1.300 ;
        RECT  0.055 0.500 0.450 0.600 ;
        RECT  0.055 1.200 0.450 1.300 ;
    END
END DEL01

MACRO DEL015
    CLASS CORE ;
    FOREIGN DEL015 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.275 2.350 1.490 ;
        RECT  2.215 0.275 2.250 0.645 ;
        RECT  2.215 1.050 2.250 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.900 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.080 0.750 2.160 0.920 ;
        RECT  1.990 0.275 2.080 0.920 ;
        RECT  1.415 0.275 1.990 0.365 ;
        RECT  1.525 0.475 1.635 1.480 ;
        RECT  1.310 0.275 1.415 1.450 ;
        RECT  1.215 0.275 1.310 0.405 ;
        RECT  1.215 1.320 1.310 1.450 ;
        RECT  1.135 0.750 1.220 0.920 ;
        RECT  1.015 0.490 1.135 1.180 ;
        RECT  0.755 0.275 0.885 1.480 ;
        RECT  0.470 0.500 0.600 1.130 ;
        RECT  0.190 0.500 0.470 0.600 ;
        RECT  0.185 1.030 0.470 1.130 ;
        RECT  0.075 0.350 0.190 0.600 ;
        RECT  0.070 1.030 0.185 1.485 ;
    END
END DEL015

MACRO DEL02
    CLASS CORE ;
    FOREIGN DEL02 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.275 2.550 1.490 ;
        RECT  2.415 0.275 2.450 0.675 ;
        RECT  2.415 1.040 2.450 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.265 -0.165 2.600 0.165 ;
        RECT  2.155 -0.165 2.265 0.630 ;
        RECT  0.395 -0.165 2.155 0.165 ;
        RECT  0.395 0.300 0.500 0.410 ;
        RECT  0.285 -0.165 0.395 0.410 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.265 1.635 2.600 1.965 ;
        RECT  2.155 1.075 2.265 1.965 ;
        RECT  0.445 1.635 2.155 1.965 ;
        RECT  0.335 1.260 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.240 0.740 2.350 0.950 ;
        RECT  2.015 0.840 2.240 0.950 ;
        RECT  1.905 0.840 2.015 1.470 ;
        RECT  1.485 1.360 1.905 1.470 ;
        RECT  1.635 0.420 1.745 1.250 ;
        RECT  1.385 0.420 1.485 1.470 ;
        RECT  1.220 0.730 1.295 0.940 ;
        RECT  1.110 0.330 1.220 1.470 ;
        RECT  0.850 0.330 0.960 1.470 ;
        RECT  0.630 0.500 0.740 1.100 ;
        RECT  0.185 0.500 0.630 0.600 ;
        RECT  0.185 1.000 0.630 1.100 ;
        RECT  0.075 0.375 0.185 0.600 ;
        RECT  0.075 1.000 0.185 1.470 ;
    END
END DEL02

MACRO DEL1
    CLASS CORE ;
    FOREIGN DEL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1310 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.280 3.350 1.490 ;
        RECT  3.215 0.280 3.250 0.490 ;
        RECT  3.215 1.280 3.250 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.940 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 -0.165 3.400 0.165 ;
        RECT  2.900 0.300 3.105 0.410 ;
        RECT  2.790 -0.165 2.900 0.410 ;
        RECT  0.610 -0.165 2.790 0.165 ;
        RECT  0.500 -0.165 0.610 0.410 ;
        RECT  0.000 -0.165 0.500 0.165 ;
        RECT  0.295 0.300 0.500 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.065 1.635 3.400 1.965 ;
        RECT  2.955 1.270 3.065 1.965 ;
        RECT  0.445 1.635 2.955 1.965 ;
        RECT  0.335 1.270 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.060 0.585 3.160 1.150 ;
        RECT  1.885 0.585 3.060 0.695 ;
        RECT  1.885 1.040 3.060 1.150 ;
        RECT  1.625 0.785 2.675 0.890 ;
        RECT  1.775 0.275 1.885 0.695 ;
        RECT  1.775 1.040 1.885 1.470 ;
        RECT  1.515 0.275 1.625 1.470 ;
        RECT  0.585 0.780 1.235 0.890 ;
        RECT  0.475 0.500 0.585 1.150 ;
        RECT  0.185 0.500 0.475 0.600 ;
        RECT  0.185 1.050 0.475 1.150 ;
        RECT  0.075 0.350 0.185 0.600 ;
        RECT  0.075 1.050 0.185 1.480 ;
    END
END DEL1

MACRO DEL2
    CLASS CORE ;
    FOREIGN DEL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.245 0.310 5.350 1.490 ;
        RECT  5.125 0.310 5.245 0.440 ;
        RECT  5.125 1.330 5.245 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.015 -0.165 5.400 0.165 ;
        RECT  4.905 -0.165 5.015 0.475 ;
        RECT  2.745 -0.165 4.905 0.165 ;
        RECT  2.615 -0.165 2.745 0.470 ;
        RECT  0.405 -0.165 2.615 0.165 ;
        RECT  0.405 0.305 0.525 0.410 ;
        RECT  0.295 -0.165 0.405 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.015 1.635 5.400 1.965 ;
        RECT  4.905 1.260 5.015 1.965 ;
        RECT  2.750 1.635 4.905 1.965 ;
        RECT  2.615 1.275 2.750 1.965 ;
        RECT  0.455 1.635 2.615 1.965 ;
        RECT  0.345 1.250 0.455 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.050 0.585 5.155 1.150 ;
        RECT  4.020 0.585 5.050 0.690 ;
        RECT  4.020 1.040 5.050 1.150 ;
        RECT  3.730 0.780 4.775 0.890 ;
        RECT  3.910 0.325 4.020 0.690 ;
        RECT  3.910 1.040 4.020 1.470 ;
        RECT  3.620 0.325 3.730 1.470 ;
        RECT  2.740 0.780 3.480 0.890 ;
        RECT  2.630 0.585 2.740 1.150 ;
        RECT  1.740 0.585 2.630 0.690 ;
        RECT  1.740 1.040 2.630 1.150 ;
        RECT  1.450 0.780 2.485 0.890 ;
        RECT  1.630 0.275 1.740 0.690 ;
        RECT  1.630 1.040 1.740 1.470 ;
        RECT  1.340 0.275 1.450 1.470 ;
        RECT  0.620 0.780 1.225 0.890 ;
        RECT  0.510 0.500 0.620 1.140 ;
        RECT  0.195 0.500 0.510 0.600 ;
        RECT  0.185 1.040 0.510 1.140 ;
        RECT  0.065 0.390 0.195 0.600 ;
        RECT  0.075 1.040 0.185 1.470 ;
    END
END DEL2

MACRO DEL3
    CLASS CORE ;
    FOREIGN DEL3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.845 0.310 5.950 1.490 ;
        RECT  5.725 0.310 5.845 0.440 ;
        RECT  5.725 1.330 5.845 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.615 -0.165 6.000 0.165 ;
        RECT  5.505 -0.165 5.615 0.475 ;
        RECT  3.035 -0.165 5.505 0.165 ;
        RECT  2.905 -0.165 3.035 0.470 ;
        RECT  0.495 -0.165 2.905 0.165 ;
        RECT  0.305 -0.165 0.495 0.410 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.615 1.635 6.000 1.965 ;
        RECT  5.505 1.260 5.615 1.965 ;
        RECT  3.040 1.635 5.505 1.965 ;
        RECT  2.905 1.275 3.040 1.965 ;
        RECT  0.445 1.635 2.905 1.965 ;
        RECT  0.335 1.250 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.650 0.585 5.755 1.150 ;
        RECT  4.455 0.585 5.650 0.690 ;
        RECT  4.455 1.040 5.650 1.150 ;
        RECT  4.185 0.780 5.370 0.890 ;
        RECT  4.345 0.325 4.455 0.690 ;
        RECT  4.345 1.040 4.455 1.470 ;
        RECT  4.075 0.325 4.185 1.470 ;
        RECT  3.030 0.780 3.910 0.890 ;
        RECT  2.920 0.585 3.030 1.150 ;
        RECT  1.865 0.585 2.920 0.690 ;
        RECT  1.865 1.040 2.920 1.150 ;
        RECT  1.595 0.780 2.780 0.890 ;
        RECT  1.755 0.275 1.865 0.690 ;
        RECT  1.755 1.040 1.865 1.470 ;
        RECT  1.485 0.275 1.595 1.470 ;
        RECT  0.600 0.780 1.375 0.890 ;
        RECT  0.490 0.500 0.600 1.140 ;
        RECT  0.195 0.500 0.490 0.600 ;
        RECT  0.185 1.040 0.490 1.140 ;
        RECT  0.065 0.390 0.195 0.600 ;
        RECT  0.075 1.040 0.185 1.470 ;
    END
END DEL3

MACRO DEL4
    CLASS CORE ;
    FOREIGN DEL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.045 0.275 6.150 1.490 ;
        RECT  5.995 0.275 6.045 0.475 ;
        RECT  6.000 1.270 6.045 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.855 -0.165 6.200 0.165 ;
        RECT  5.715 -0.165 5.855 0.475 ;
        RECT  3.135 -0.165 5.715 0.165 ;
        RECT  3.005 -0.165 3.135 0.470 ;
        RECT  0.495 -0.165 3.005 0.165 ;
        RECT  0.295 -0.165 0.495 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.835 1.635 6.200 1.965 ;
        RECT  5.725 1.260 5.835 1.965 ;
        RECT  3.140 1.635 5.725 1.965 ;
        RECT  3.005 1.275 3.140 1.965 ;
        RECT  0.445 1.635 3.005 1.965 ;
        RECT  0.335 1.250 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.865 0.585 5.955 1.150 ;
        RECT  4.605 0.585 5.865 0.690 ;
        RECT  4.605 1.040 5.865 1.150 ;
        RECT  4.325 0.780 5.530 0.890 ;
        RECT  4.495 0.325 4.605 0.690 ;
        RECT  4.495 1.040 4.605 1.470 ;
        RECT  4.215 0.325 4.325 1.470 ;
        RECT  3.205 0.780 4.050 0.890 ;
        RECT  3.095 0.585 3.205 1.150 ;
        RECT  1.925 0.585 3.095 0.690 ;
        RECT  1.925 1.040 3.095 1.150 ;
        RECT  1.645 0.780 2.880 0.890 ;
        RECT  1.815 0.325 1.925 0.690 ;
        RECT  1.815 1.040 1.925 1.470 ;
        RECT  1.535 0.325 1.645 1.470 ;
        RECT  0.600 0.780 1.395 0.890 ;
        RECT  0.490 0.500 0.600 1.140 ;
        RECT  0.195 0.500 0.490 0.600 ;
        RECT  0.185 1.040 0.490 1.140 ;
        RECT  0.065 0.390 0.195 0.600 ;
        RECT  0.075 1.040 0.185 1.470 ;
    END
END DEL4

MACRO DFCND1
    CLASS CORE ;
    FOREIGN DFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.285 4.755 1.490 ;
        RECT  4.625 0.285 4.650 0.675 ;
        RECT  4.625 1.040 4.650 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1430 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.305 4.355 1.125 ;
        RECT  4.065 0.305 4.245 0.415 ;
        RECT  4.075 1.030 4.245 1.125 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0486 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.255 0.910 ;
        RECT  1.050 0.730 1.155 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.650 0.155 1.110 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.490 3.755 0.890 ;
        RECT  3.445 0.710 3.650 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 -0.165 4.800 0.165 ;
        RECT  3.390 -0.165 3.560 0.590 ;
        RECT  2.045 -0.165 3.390 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.895 -0.165 1.915 0.165 ;
        RECT  0.705 -0.165 0.895 0.355 ;
        RECT  0.000 -0.165 0.705 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.635 4.800 1.965 ;
        RECT  0.340 1.475 0.510 1.965 ;
        RECT  0.000 1.635 0.340 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.535 0.775 4.560 0.945 ;
        RECT  4.445 0.775 4.535 1.315 ;
        RECT  3.160 1.225 4.445 1.315 ;
        RECT  3.990 0.780 4.135 0.890 ;
        RECT  3.960 0.505 3.990 0.890 ;
        RECT  3.855 0.505 3.960 1.135 ;
        RECT  3.350 1.025 3.855 1.135 ;
        RECT  3.630 1.435 3.855 1.525 ;
        RECT  3.540 1.405 3.630 1.525 ;
        RECT  2.960 1.405 3.540 1.495 ;
        RECT  3.250 0.735 3.350 1.135 ;
        RECT  3.100 0.525 3.300 0.625 ;
        RECT  3.225 0.735 3.250 0.945 ;
        RECT  3.100 1.035 3.160 1.315 ;
        RECT  2.890 0.275 3.120 0.435 ;
        RECT  3.050 0.525 3.100 1.315 ;
        RECT  3.010 0.525 3.050 1.125 ;
        RECT  2.800 0.665 3.010 0.775 ;
        RECT  2.900 1.215 2.960 1.495 ;
        RECT  2.860 0.945 2.900 1.495 ;
        RECT  2.225 0.275 2.890 0.365 ;
        RECT  2.790 0.945 2.860 1.320 ;
        RECT  2.675 0.945 2.790 1.045 ;
        RECT  2.600 1.410 2.770 1.520 ;
        RECT  2.425 1.175 2.685 1.280 ;
        RECT  2.565 0.455 2.675 1.045 ;
        RECT  0.720 1.430 2.600 1.520 ;
        RECT  2.315 0.455 2.425 1.280 ;
        RECT  1.705 1.010 2.315 1.110 ;
        RECT  2.135 0.275 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.470 1.210 2.135 1.340 ;
        RECT  1.455 0.720 2.095 0.820 ;
        RECT  1.595 0.910 1.705 1.110 ;
        RECT  1.570 0.275 1.660 0.605 ;
        RECT  1.105 0.275 1.570 0.365 ;
        RECT  1.380 0.505 1.455 1.110 ;
        RECT  1.355 0.505 1.380 1.320 ;
        RECT  1.200 0.505 1.355 0.615 ;
        RECT  1.270 1.020 1.355 1.320 ;
        RECT  1.200 1.200 1.270 1.320 ;
        RECT  1.005 0.275 1.105 0.580 ;
        RECT  0.685 0.470 1.005 0.580 ;
        RECT  0.685 0.790 0.830 0.900 ;
        RECT  0.620 1.265 0.720 1.520 ;
        RECT  0.575 0.470 0.685 1.175 ;
        RECT  0.410 1.265 0.620 1.365 ;
        RECT  0.310 0.440 0.410 1.365 ;
        RECT  0.180 0.440 0.310 0.540 ;
        RECT  0.185 1.255 0.310 1.365 ;
        RECT  0.075 1.255 0.185 1.445 ;
        RECT  0.080 0.350 0.180 0.540 ;
    END
END DFCND1

MACRO DFCND2
    CLASS CORE ;
    FOREIGN DFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.150 1.090 5.310 1.220 ;
        RECT  5.150 0.285 5.260 0.690 ;
        RECT  5.050 0.580 5.150 1.220 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.580 4.950 1.220 ;
        RECT  4.760 0.580 4.850 0.690 ;
        RECT  4.600 1.090 4.850 1.220 ;
        RECT  4.650 0.285 4.760 0.690 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0486 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.255 0.910 ;
        RECT  1.050 0.730 1.155 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.650 0.155 1.110 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0934 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.490 3.755 0.890 ;
        RECT  3.445 0.710 3.650 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 -0.165 5.600 0.165 ;
        RECT  5.410 -0.165 5.520 0.685 ;
        RECT  4.505 -0.165 5.410 0.165 ;
        RECT  4.335 -0.165 4.505 0.585 ;
        RECT  3.560 -0.165 4.335 0.165 ;
        RECT  3.390 -0.165 3.560 0.590 ;
        RECT  2.045 -0.165 3.390 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.895 -0.165 1.915 0.165 ;
        RECT  0.705 -0.165 0.895 0.355 ;
        RECT  0.000 -0.165 0.705 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.635 5.600 1.965 ;
        RECT  0.340 1.475 0.510 1.965 ;
        RECT  0.000 1.635 0.340 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.420 0.790 5.510 1.430 ;
        RECT  5.260 0.790 5.420 0.900 ;
        RECT  4.095 1.340 5.420 1.430 ;
        RECT  3.990 0.780 4.740 0.890 ;
        RECT  3.990 1.025 4.310 1.135 ;
        RECT  3.975 1.225 4.095 1.430 ;
        RECT  3.880 0.505 3.990 1.135 ;
        RECT  3.160 1.225 3.975 1.315 ;
        RECT  3.350 1.025 3.880 1.135 ;
        RECT  3.630 1.435 3.855 1.525 ;
        RECT  3.540 1.405 3.630 1.525 ;
        RECT  2.960 1.405 3.540 1.495 ;
        RECT  3.250 0.735 3.350 1.135 ;
        RECT  3.100 0.525 3.300 0.625 ;
        RECT  3.225 0.735 3.250 0.945 ;
        RECT  3.100 1.035 3.160 1.315 ;
        RECT  2.890 0.275 3.120 0.435 ;
        RECT  3.050 0.525 3.100 1.315 ;
        RECT  3.010 0.525 3.050 1.125 ;
        RECT  2.800 0.665 3.010 0.775 ;
        RECT  2.900 1.215 2.960 1.495 ;
        RECT  2.860 0.945 2.900 1.495 ;
        RECT  2.225 0.275 2.890 0.365 ;
        RECT  2.790 0.945 2.860 1.320 ;
        RECT  2.675 0.945 2.790 1.045 ;
        RECT  2.600 1.410 2.770 1.520 ;
        RECT  2.425 1.175 2.685 1.280 ;
        RECT  2.565 0.455 2.675 1.045 ;
        RECT  0.720 1.430 2.600 1.520 ;
        RECT  2.315 0.455 2.425 1.280 ;
        RECT  1.705 1.010 2.315 1.110 ;
        RECT  2.135 0.275 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.470 1.210 2.135 1.340 ;
        RECT  1.455 0.720 2.095 0.820 ;
        RECT  1.595 0.910 1.705 1.110 ;
        RECT  1.570 0.275 1.660 0.605 ;
        RECT  1.105 0.275 1.570 0.365 ;
        RECT  1.380 0.505 1.455 1.110 ;
        RECT  1.355 0.505 1.380 1.320 ;
        RECT  1.200 0.505 1.355 0.615 ;
        RECT  1.270 1.020 1.355 1.320 ;
        RECT  1.200 1.200 1.270 1.320 ;
        RECT  1.005 0.275 1.105 0.600 ;
        RECT  0.685 0.490 1.005 0.600 ;
        RECT  0.685 0.790 0.830 0.900 ;
        RECT  0.620 1.265 0.720 1.520 ;
        RECT  0.575 0.490 0.685 1.175 ;
        RECT  0.410 1.265 0.620 1.365 ;
        RECT  0.310 0.440 0.410 1.365 ;
        RECT  0.180 0.440 0.310 0.540 ;
        RECT  0.185 1.255 0.310 1.365 ;
        RECT  0.075 1.255 0.185 1.445 ;
        RECT  0.080 0.350 0.180 0.540 ;
    END
END DFCND2

MACRO DFCND4
    CLASS CORE ;
    FOREIGN DFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.150 0.285 6.260 1.500 ;
        RECT  5.950 0.505 6.150 1.210 ;
        RECT  5.760 0.505 5.950 0.675 ;
        RECT  5.760 1.040 5.950 1.210 ;
        RECT  5.650 0.285 5.760 0.675 ;
        RECT  5.650 1.040 5.760 1.500 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 1.050 5.310 1.220 ;
        RECT  5.150 0.285 5.260 0.675 ;
        RECT  5.050 0.505 5.150 0.675 ;
        RECT  4.760 0.505 5.050 1.220 ;
        RECT  4.750 0.285 4.760 1.220 ;
        RECT  4.650 0.285 4.750 0.675 ;
        RECT  4.600 1.050 4.750 1.220 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0486 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.710 1.255 0.910 ;
        RECT  1.050 0.710 1.155 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.650 0.155 1.110 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0933 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.490 3.755 0.890 ;
        RECT  3.445 0.710 3.650 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.520 -0.165 6.600 0.165 ;
        RECT  6.410 -0.165 6.520 0.695 ;
        RECT  4.485 -0.165 6.410 0.165 ;
        RECT  4.355 -0.165 4.485 0.675 ;
        RECT  3.560 -0.165 4.355 0.165 ;
        RECT  3.390 -0.165 3.560 0.590 ;
        RECT  2.045 -0.165 3.390 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.930 -0.165 1.915 0.165 ;
        RECT  0.760 -0.165 0.930 0.440 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.520 1.635 6.600 1.965 ;
        RECT  6.410 1.040 6.520 1.965 ;
        RECT  0.000 1.635 6.410 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.760 0.505 5.850 0.675 ;
        RECT  5.760 1.040 5.850 1.210 ;
        RECT  5.650 0.285 5.760 0.675 ;
        RECT  5.650 1.040 5.760 1.500 ;
        RECT  5.150 1.050 5.310 1.220 ;
        RECT  5.150 0.285 5.260 0.675 ;
        RECT  4.600 1.050 4.650 1.220 ;
        RECT  5.520 0.780 5.755 0.890 ;
        RECT  5.430 0.780 5.520 1.430 ;
        RECT  4.095 1.340 5.430 1.430 ;
        RECT  3.990 0.780 4.655 0.890 ;
        RECT  3.990 1.025 4.310 1.135 ;
        RECT  3.975 1.225 4.095 1.430 ;
        RECT  3.880 0.490 3.990 1.135 ;
        RECT  3.160 1.225 3.975 1.315 ;
        RECT  3.350 1.025 3.880 1.135 ;
        RECT  3.630 1.435 3.855 1.525 ;
        RECT  3.540 1.405 3.630 1.525 ;
        RECT  2.960 1.405 3.540 1.495 ;
        RECT  3.250 0.735 3.350 1.135 ;
        RECT  3.100 0.525 3.300 0.625 ;
        RECT  3.225 0.735 3.250 0.945 ;
        RECT  3.100 1.035 3.160 1.315 ;
        RECT  2.890 0.275 3.120 0.435 ;
        RECT  3.050 0.525 3.100 1.315 ;
        RECT  3.010 0.525 3.050 1.125 ;
        RECT  2.800 0.665 3.010 0.775 ;
        RECT  2.900 1.215 2.960 1.495 ;
        RECT  2.860 0.945 2.900 1.495 ;
        RECT  2.225 0.275 2.890 0.365 ;
        RECT  2.790 0.945 2.860 1.320 ;
        RECT  2.675 0.945 2.790 1.045 ;
        RECT  2.600 1.410 2.770 1.525 ;
        RECT  2.425 1.175 2.685 1.280 ;
        RECT  2.565 0.455 2.675 1.045 ;
        RECT  0.410 1.430 2.600 1.525 ;
        RECT  2.315 0.455 2.425 1.280 ;
        RECT  1.705 1.010 2.315 1.110 ;
        RECT  2.135 0.275 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.470 1.210 2.135 1.340 ;
        RECT  1.455 0.720 2.095 0.820 ;
        RECT  1.595 0.910 1.705 1.110 ;
        RECT  1.570 0.275 1.660 0.605 ;
        RECT  1.120 0.275 1.570 0.365 ;
        RECT  1.380 0.505 1.455 1.110 ;
        RECT  1.355 0.505 1.380 1.320 ;
        RECT  1.210 0.505 1.355 0.615 ;
        RECT  1.270 1.020 1.355 1.320 ;
        RECT  1.200 1.200 1.270 1.320 ;
        RECT  1.030 0.275 1.120 0.620 ;
        RECT  0.795 0.530 1.030 0.620 ;
        RECT  0.680 0.530 0.795 1.245 ;
        RECT  0.545 0.530 0.680 0.655 ;
        RECT  0.525 1.115 0.680 1.245 ;
        RECT  0.410 0.770 0.520 0.940 ;
        RECT  0.310 0.440 0.410 1.525 ;
        RECT  0.180 0.440 0.310 0.540 ;
        RECT  0.185 1.415 0.310 1.525 ;
        RECT  0.075 1.255 0.185 1.525 ;
        RECT  0.080 0.350 0.180 0.540 ;
    END
END DFCND4

MACRO DFCNQD1
    CLASS CORE ;
    FOREIGN DFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.285 4.355 1.490 ;
        RECT  4.215 0.285 4.250 0.675 ;
        RECT  4.215 1.040 4.250 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0486 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.255 0.910 ;
        RECT  1.045 0.730 1.155 1.320 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.710 0.200 0.960 ;
        RECT  0.045 0.710 0.155 1.090 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0665 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.550 1.090 ;
        RECT  3.410 0.895 3.450 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.430 -0.165 4.400 0.165 ;
        RECT  3.260 -0.165 3.430 0.420 ;
        RECT  2.045 -0.165 3.260 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.875 -0.165 1.915 0.165 ;
        RECT  0.765 -0.165 0.875 0.415 ;
        RECT  0.000 -0.165 0.765 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.400 1.635 4.400 1.965 ;
        RECT  3.260 1.365 3.400 1.965 ;
        RECT  0.000 1.635 3.260 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.070 0.780 4.160 0.890 ;
        RECT  3.960 0.510 4.070 1.470 ;
        RECT  3.270 0.510 3.960 0.620 ;
        RECT  3.525 1.365 3.960 1.470 ;
        RECT  3.740 0.750 3.850 1.275 ;
        RECT  2.900 1.180 3.740 1.275 ;
        RECT  3.160 0.510 3.270 1.085 ;
        RECT  2.910 0.325 3.020 0.925 ;
        RECT  2.225 0.325 2.910 0.415 ;
        RECT  2.790 1.035 2.900 1.275 ;
        RECT  2.675 1.035 2.790 1.125 ;
        RECT  2.600 1.410 2.770 1.525 ;
        RECT  2.425 1.215 2.680 1.310 ;
        RECT  2.565 0.505 2.675 1.125 ;
        RECT  0.410 1.435 2.600 1.525 ;
        RECT  2.315 0.505 2.425 1.310 ;
        RECT  1.705 1.010 2.315 1.110 ;
        RECT  2.135 0.325 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.465 1.210 2.135 1.345 ;
        RECT  1.455 0.720 2.095 0.820 ;
        RECT  1.595 0.910 1.705 1.110 ;
        RECT  1.570 0.275 1.660 0.605 ;
        RECT  1.105 0.275 1.570 0.375 ;
        RECT  1.355 0.505 1.455 1.110 ;
        RECT  1.200 0.505 1.355 0.615 ;
        RECT  1.245 1.020 1.355 1.340 ;
        RECT  1.005 0.275 1.105 0.625 ;
        RECT  0.685 0.535 1.005 0.625 ;
        RECT  0.685 0.835 0.830 0.945 ;
        RECT  0.575 0.495 0.685 1.325 ;
        RECT  0.310 0.490 0.410 1.525 ;
        RECT  0.045 0.490 0.310 0.600 ;
        RECT  0.045 1.200 0.310 1.310 ;
    END
END DFCNQD1

MACRO DFCNQD2
    CLASS CORE ;
    FOREIGN DFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.575 4.750 1.490 ;
        RECT  4.640 0.575 4.650 0.675 ;
        RECT  4.565 1.040 4.650 1.490 ;
        RECT  4.530 0.285 4.640 0.675 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0486 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.255 0.910 ;
        RECT  1.045 0.730 1.155 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.650 0.155 1.110 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0963 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.550 1.090 ;
        RECT  3.420 0.710 3.450 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.420 -0.165 5.000 0.165 ;
        RECT  3.250 -0.165 3.420 0.420 ;
        RECT  2.045 -0.165 3.250 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.875 -0.165 1.915 0.165 ;
        RECT  0.765 -0.165 0.875 0.445 ;
        RECT  0.000 -0.165 0.765 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.405 1.635 5.000 1.965 ;
        RECT  3.250 1.380 3.405 1.965 ;
        RECT  0.000 1.635 3.250 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.420 0.765 4.540 0.935 ;
        RECT  4.310 0.510 4.420 1.470 ;
        RECT  3.270 0.510 4.310 0.620 ;
        RECT  3.515 1.360 4.310 1.470 ;
        RECT  3.825 0.730 3.935 1.270 ;
        RECT  2.900 1.180 3.825 1.270 ;
        RECT  3.160 0.510 3.270 0.940 ;
        RECT  2.910 0.325 3.020 0.925 ;
        RECT  2.225 0.325 2.910 0.415 ;
        RECT  2.790 1.035 2.900 1.270 ;
        RECT  2.675 1.035 2.790 1.125 ;
        RECT  0.410 1.435 2.790 1.525 ;
        RECT  2.425 1.215 2.680 1.325 ;
        RECT  2.565 0.505 2.675 1.125 ;
        RECT  2.315 0.505 2.425 1.325 ;
        RECT  1.705 1.010 2.315 1.110 ;
        RECT  2.135 0.325 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.890 1.255 2.135 1.345 ;
        RECT  1.455 0.720 2.095 0.820 ;
        RECT  1.770 1.210 1.890 1.345 ;
        RECT  1.465 1.210 1.770 1.310 ;
        RECT  1.595 0.910 1.705 1.110 ;
        RECT  1.570 0.275 1.660 0.605 ;
        RECT  1.105 0.275 1.570 0.365 ;
        RECT  1.355 0.505 1.455 1.110 ;
        RECT  1.200 0.505 1.355 0.615 ;
        RECT  1.245 1.020 1.355 1.340 ;
        RECT  1.005 0.275 1.105 0.625 ;
        RECT  0.685 0.535 1.005 0.625 ;
        RECT  0.685 0.790 0.830 0.900 ;
        RECT  0.575 0.495 0.685 1.325 ;
        RECT  0.310 0.440 0.410 1.525 ;
        RECT  0.180 0.440 0.310 0.540 ;
        RECT  0.075 1.255 0.310 1.445 ;
        RECT  0.080 0.350 0.180 0.540 ;
    END
END DFCNQD2

MACRO DFCNQD4
    CLASS CORE ;
    FOREIGN DFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.150 0.275 5.260 0.675 ;
        RECT  5.150 1.040 5.260 1.500 ;
        RECT  5.050 0.505 5.150 0.675 ;
        RECT  5.050 1.040 5.150 1.210 ;
        RECT  4.760 0.505 5.050 1.210 ;
        RECT  4.750 0.275 4.760 1.500 ;
        RECT  4.650 0.275 4.750 0.675 ;
        RECT  4.650 1.040 4.750 1.500 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0486 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.255 0.910 ;
        RECT  1.045 0.730 1.155 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.700 0.200 0.940 ;
        RECT  0.045 0.700 0.155 1.110 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0981 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.490 3.755 0.890 ;
        RECT  3.445 0.710 3.650 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 -0.165 5.600 0.165 ;
        RECT  5.410 -0.165 5.520 0.695 ;
        RECT  4.475 -0.165 5.410 0.165 ;
        RECT  4.365 -0.165 4.475 0.670 ;
        RECT  3.560 -0.165 4.365 0.165 ;
        RECT  3.390 -0.165 3.560 0.620 ;
        RECT  2.045 -0.165 3.390 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.895 -0.165 1.915 0.165 ;
        RECT  0.790 -0.165 0.895 0.445 ;
        RECT  0.000 -0.165 0.790 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.635 5.600 1.965 ;
        RECT  5.410 1.040 5.520 1.965 ;
        RECT  3.425 1.635 5.410 1.965 ;
        RECT  3.285 1.455 3.425 1.965 ;
        RECT  0.000 1.635 3.285 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.150 0.275 5.260 0.675 ;
        RECT  5.150 1.040 5.260 1.500 ;
        RECT  4.260 0.780 4.655 0.890 ;
        RECT  4.150 0.490 4.260 1.500 ;
        RECT  3.845 0.490 4.150 0.600 ;
        RECT  3.350 1.025 4.150 1.135 ;
        RECT  3.625 1.425 3.855 1.525 ;
        RECT  3.535 1.245 3.625 1.525 ;
        RECT  2.900 1.245 3.535 1.335 ;
        RECT  3.250 0.735 3.350 1.135 ;
        RECT  2.960 0.525 3.300 0.625 ;
        RECT  3.225 0.735 3.250 0.945 ;
        RECT  2.890 0.275 3.120 0.435 ;
        RECT  2.850 0.525 2.960 0.825 ;
        RECT  2.790 0.945 2.900 1.335 ;
        RECT  2.225 0.275 2.890 0.365 ;
        RECT  2.675 0.945 2.790 1.045 ;
        RECT  2.600 1.430 2.770 1.545 ;
        RECT  2.425 1.175 2.685 1.280 ;
        RECT  2.565 0.455 2.675 1.045 ;
        RECT  0.410 1.430 2.600 1.520 ;
        RECT  2.315 0.455 2.425 1.280 ;
        RECT  1.705 1.010 2.315 1.110 ;
        RECT  2.135 0.275 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.465 1.210 2.135 1.340 ;
        RECT  1.455 0.720 2.095 0.820 ;
        RECT  1.595 0.910 1.705 1.110 ;
        RECT  1.570 0.275 1.660 0.605 ;
        RECT  1.105 0.275 1.570 0.365 ;
        RECT  1.355 0.505 1.455 1.110 ;
        RECT  1.200 0.505 1.355 0.615 ;
        RECT  1.245 1.020 1.355 1.340 ;
        RECT  1.005 0.275 1.105 0.630 ;
        RECT  0.790 0.535 1.005 0.630 ;
        RECT  0.680 0.535 0.790 1.320 ;
        RECT  0.525 0.535 0.680 0.655 ;
        RECT  0.525 1.210 0.680 1.320 ;
        RECT  0.410 0.750 0.520 0.920 ;
        RECT  0.310 0.440 0.410 1.520 ;
        RECT  0.180 0.440 0.310 0.540 ;
        RECT  0.045 1.220 0.310 1.330 ;
        RECT  0.080 0.350 0.180 0.540 ;
    END
END DFCNQD4

MACRO DFCSND1
    CLASS CORE ;
    FOREIGN DFCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0755 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.275 5.550 1.490 ;
        RECT  5.420 0.275 5.450 0.675 ;
        RECT  5.420 1.045 5.450 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.455 5.150 1.175 ;
        RECT  4.870 0.455 5.050 0.625 ;
        RECT  4.985 1.065 5.050 1.175 ;
        RECT  4.850 1.065 4.985 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0533 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.760 1.290 0.945 ;
        RECT  1.150 0.800 1.180 0.945 ;
        RECT  1.050 0.800 1.150 1.300 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0737 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.710 4.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.220 -0.165 5.600 0.165 ;
        RECT  4.045 -0.165 4.220 0.420 ;
        RECT  2.220 -0.165 4.045 0.165 ;
        RECT  2.050 -0.165 2.220 0.355 ;
        RECT  0.945 -0.165 2.050 0.165 ;
        RECT  0.835 -0.165 0.945 0.480 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.260 1.635 5.600 1.965 ;
        RECT  5.130 1.320 5.260 1.965 ;
        RECT  3.650 1.635 5.130 1.965 ;
        RECT  3.485 1.435 3.650 1.965 ;
        RECT  3.480 1.435 3.485 1.525 ;
        RECT  2.760 1.635 3.485 1.965 ;
        RECT  2.570 1.425 2.760 1.965 ;
        RECT  0.000 1.635 2.570 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.330 0.750 5.360 0.920 ;
        RECT  5.240 0.275 5.330 0.920 ;
        RECT  4.445 0.275 5.240 0.365 ;
        RECT  4.760 0.730 4.910 0.945 ;
        RECT  4.655 0.455 4.760 1.500 ;
        RECT  4.550 0.455 4.655 0.580 ;
        RECT  4.090 1.390 4.655 1.500 ;
        RECT  4.445 0.765 4.555 1.295 ;
        RECT  4.355 0.275 4.445 0.620 ;
        RECT  3.870 1.205 4.445 1.295 ;
        RECT  3.360 0.510 4.355 0.620 ;
        RECT  4.000 1.390 4.090 1.545 ;
        RECT  3.830 1.435 4.000 1.545 ;
        RECT  3.625 1.025 3.955 1.115 ;
        RECT  3.780 1.205 3.870 1.335 ;
        RECT  3.175 1.245 3.780 1.335 ;
        RECT  3.360 1.025 3.625 1.155 ;
        RECT  3.270 0.510 3.360 1.155 ;
        RECT  2.435 0.315 3.350 0.415 ;
        RECT  3.055 0.570 3.270 0.695 ;
        RECT  3.070 0.825 3.175 1.335 ;
        RECT  2.945 0.825 3.070 0.915 ;
        RECT  2.885 1.245 2.975 1.525 ;
        RECT  2.835 0.525 2.945 0.915 ;
        RECT  2.680 1.055 2.940 1.155 ;
        RECT  2.415 1.245 2.885 1.335 ;
        RECT  2.560 0.505 2.680 1.155 ;
        RECT  2.105 1.055 2.560 1.155 ;
        RECT  2.345 0.315 2.435 0.535 ;
        RECT  2.325 1.245 2.415 1.525 ;
        RECT  1.920 0.445 2.345 0.535 ;
        RECT  1.555 1.425 2.325 1.525 ;
        RECT  2.200 0.625 2.315 0.940 ;
        RECT  1.510 0.625 2.200 0.715 ;
        RECT  2.015 0.805 2.105 1.155 ;
        RECT  1.630 0.805 2.015 0.895 ;
        RECT  1.835 1.005 1.925 1.325 ;
        RECT  1.830 0.275 1.920 0.535 ;
        RECT  1.460 1.235 1.835 1.325 ;
        RECT  1.155 0.275 1.830 0.375 ;
        RECT  1.345 1.425 1.555 1.545 ;
        RECT  1.505 0.545 1.510 0.715 ;
        RECT  1.415 0.545 1.505 1.145 ;
        RECT  1.285 0.545 1.415 0.650 ;
        RECT  1.350 1.055 1.415 1.145 ;
        RECT  1.260 1.055 1.350 1.335 ;
        RECT  0.450 1.425 1.345 1.525 ;
        RECT  1.065 0.275 1.155 0.660 ;
        RECT  0.800 0.570 1.065 0.660 ;
        RECT  0.685 0.570 0.800 1.315 ;
        RECT  0.660 0.355 0.685 1.315 ;
        RECT  0.575 0.355 0.660 0.660 ;
        RECT  0.540 1.205 0.660 1.315 ;
        RECT  0.450 0.750 0.520 0.920 ;
        RECT  0.360 0.505 0.450 1.525 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.435 0.360 1.525 ;
        RECT  0.075 0.365 0.185 0.595 ;
        RECT  0.075 1.205 0.185 1.525 ;
    END
END DFCSND1

MACRO DFCSND2
    CLASS CORE ;
    FOREIGN DFCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0755 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.600 6.150 1.145 ;
        RECT  5.950 0.600 6.050 0.690 ;
        RECT  5.950 1.045 6.050 1.145 ;
        RECT  5.765 0.275 5.950 0.690 ;
        RECT  5.765 1.045 5.950 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 1.110 5.550 1.490 ;
        RECT  5.375 0.475 5.475 1.490 ;
        RECT  5.275 0.475 5.375 0.660 ;
        RECT  5.275 1.080 5.375 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0533 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.760 1.290 0.945 ;
        RECT  1.150 0.800 1.180 0.945 ;
        RECT  1.050 0.800 1.150 1.300 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1289 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.900 0.635 5.005 0.940 ;
        RECT  4.550 0.635 4.900 0.725 ;
        RECT  4.450 0.635 4.550 1.100 ;
        RECT  4.440 0.780 4.450 1.100 ;
        RECT  4.125 0.780 4.440 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.160 -0.165 6.200 0.165 ;
        RECT  3.985 -0.165 4.160 0.420 ;
        RECT  2.220 -0.165 3.985 0.165 ;
        RECT  2.050 -0.165 2.220 0.355 ;
        RECT  0.945 -0.165 2.050 0.165 ;
        RECT  0.835 -0.165 0.945 0.480 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.615 1.635 6.200 1.965 ;
        RECT  3.445 1.435 3.615 1.965 ;
        RECT  2.745 1.635 3.445 1.965 ;
        RECT  2.555 1.435 2.745 1.965 ;
        RECT  0.000 1.635 2.555 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.675 0.780 5.900 0.890 ;
        RECT  5.585 0.275 5.675 0.890 ;
        RECT  4.340 0.275 5.585 0.365 ;
        RECT  5.185 0.750 5.285 0.920 ;
        RECT  5.095 0.455 5.185 1.500 ;
        RECT  4.505 0.455 5.095 0.545 ;
        RECT  4.055 1.390 5.095 1.500 ;
        RECT  4.640 0.815 4.810 1.295 ;
        RECT  3.835 1.205 4.640 1.295 ;
        RECT  4.250 0.275 4.340 0.620 ;
        RECT  3.335 0.510 4.250 0.620 ;
        RECT  3.965 1.390 4.055 1.545 ;
        RECT  3.810 1.435 3.965 1.545 ;
        RECT  3.455 1.015 3.920 1.115 ;
        RECT  3.745 1.205 3.835 1.345 ;
        RECT  3.145 1.255 3.745 1.345 ;
        RECT  3.335 1.015 3.455 1.165 ;
        RECT  2.435 0.315 3.385 0.415 ;
        RECT  3.245 0.510 3.335 1.165 ;
        RECT  3.055 0.585 3.245 0.695 ;
        RECT  3.045 0.825 3.145 1.345 ;
        RECT  2.945 0.825 3.045 0.915 ;
        RECT  2.840 1.255 2.950 1.525 ;
        RECT  2.835 0.525 2.945 0.915 ;
        RECT  2.675 1.055 2.935 1.165 ;
        RECT  2.415 1.255 2.840 1.345 ;
        RECT  2.565 0.505 2.675 1.165 ;
        RECT  2.105 1.055 2.565 1.165 ;
        RECT  2.345 0.315 2.435 0.535 ;
        RECT  2.325 1.255 2.415 1.525 ;
        RECT  1.920 0.445 2.345 0.535 ;
        RECT  1.555 1.425 2.325 1.525 ;
        RECT  2.200 0.625 2.315 0.940 ;
        RECT  1.510 0.625 2.200 0.715 ;
        RECT  2.015 0.805 2.105 1.165 ;
        RECT  1.630 0.805 2.015 0.895 ;
        RECT  1.835 1.005 1.925 1.325 ;
        RECT  1.830 0.275 1.920 0.535 ;
        RECT  1.460 1.235 1.835 1.325 ;
        RECT  1.155 0.275 1.830 0.375 ;
        RECT  1.345 1.425 1.555 1.545 ;
        RECT  1.505 0.545 1.510 0.715 ;
        RECT  1.415 0.545 1.505 1.145 ;
        RECT  1.285 0.545 1.415 0.650 ;
        RECT  1.350 1.055 1.415 1.145 ;
        RECT  1.260 1.055 1.350 1.335 ;
        RECT  0.450 1.425 1.345 1.525 ;
        RECT  1.065 0.275 1.155 0.660 ;
        RECT  0.780 0.570 1.065 0.660 ;
        RECT  0.685 0.570 0.780 1.315 ;
        RECT  0.670 0.355 0.685 1.315 ;
        RECT  0.575 0.355 0.670 0.660 ;
        RECT  0.540 1.205 0.670 1.315 ;
        RECT  0.450 0.750 0.520 0.920 ;
        RECT  0.360 0.505 0.450 1.525 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.435 0.360 1.525 ;
        RECT  0.075 0.365 0.185 0.595 ;
        RECT  0.075 1.205 0.185 1.525 ;
    END
END DFCSND2

MACRO DFCSND4
    CLASS CORE ;
    FOREIGN DFCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0755 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.325 6.950 0.635 ;
        RECT  6.850 1.100 6.950 1.410 ;
        RECT  6.550 0.325 6.850 1.410 ;
        RECT  6.235 0.325 6.550 0.635 ;
        RECT  6.235 1.100 6.550 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.510 5.925 0.690 ;
        RECT  5.850 1.310 5.925 1.490 ;
        RECT  5.550 0.510 5.850 1.490 ;
        RECT  5.275 0.510 5.550 0.690 ;
        RECT  5.235 1.310 5.550 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0533 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.760 1.290 0.945 ;
        RECT  1.150 0.800 1.180 0.945 ;
        RECT  1.050 0.800 1.150 1.300 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1289 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.900 0.635 5.005 0.920 ;
        RECT  4.550 0.635 4.900 0.725 ;
        RECT  4.450 0.635 4.550 1.100 ;
        RECT  4.440 0.780 4.450 1.100 ;
        RECT  4.125 0.780 4.440 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.160 -0.165 7.200 0.165 ;
        RECT  3.985 -0.165 4.160 0.420 ;
        RECT  2.220 -0.165 3.985 0.165 ;
        RECT  2.050 -0.165 2.220 0.355 ;
        RECT  0.945 -0.165 2.050 0.165 ;
        RECT  0.835 -0.165 0.945 0.480 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.615 1.635 7.200 1.965 ;
        RECT  3.445 1.435 3.615 1.965 ;
        RECT  2.745 1.635 3.445 1.965 ;
        RECT  2.555 1.435 2.745 1.965 ;
        RECT  0.000 1.635 2.555 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.235 0.325 6.450 0.635 ;
        RECT  6.235 1.100 6.450 1.410 ;
        RECT  5.275 0.510 5.450 0.690 ;
        RECT  5.235 1.310 5.450 1.490 ;
        RECT  6.125 0.780 6.400 0.890 ;
        RECT  6.035 0.275 6.125 0.890 ;
        RECT  4.340 0.275 6.035 0.365 ;
        RECT  5.185 0.780 5.365 0.890 ;
        RECT  5.125 0.455 5.185 1.200 ;
        RECT  5.095 0.455 5.125 1.500 ;
        RECT  4.505 0.455 5.095 0.545 ;
        RECT  5.035 1.110 5.095 1.500 ;
        RECT  4.055 1.390 5.035 1.500 ;
        RECT  4.640 0.815 4.810 1.295 ;
        RECT  3.835 1.205 4.640 1.295 ;
        RECT  4.250 0.275 4.340 0.620 ;
        RECT  3.335 0.510 4.250 0.620 ;
        RECT  3.965 1.390 4.055 1.545 ;
        RECT  3.810 1.435 3.965 1.545 ;
        RECT  3.455 1.015 3.920 1.115 ;
        RECT  3.745 1.205 3.835 1.345 ;
        RECT  3.145 1.255 3.745 1.345 ;
        RECT  3.335 1.015 3.455 1.165 ;
        RECT  2.435 0.315 3.385 0.415 ;
        RECT  3.245 0.510 3.335 1.165 ;
        RECT  3.055 0.585 3.245 0.695 ;
        RECT  3.045 0.825 3.145 1.345 ;
        RECT  2.945 0.825 3.045 0.915 ;
        RECT  2.840 1.255 2.950 1.525 ;
        RECT  2.835 0.525 2.945 0.915 ;
        RECT  2.675 1.055 2.935 1.165 ;
        RECT  2.415 1.255 2.840 1.345 ;
        RECT  2.565 0.505 2.675 1.165 ;
        RECT  2.105 1.055 2.565 1.165 ;
        RECT  2.345 0.315 2.435 0.535 ;
        RECT  2.325 1.255 2.415 1.525 ;
        RECT  1.920 0.445 2.345 0.535 ;
        RECT  1.555 1.425 2.325 1.525 ;
        RECT  2.200 0.625 2.315 0.940 ;
        RECT  1.510 0.625 2.200 0.715 ;
        RECT  2.015 0.805 2.105 1.165 ;
        RECT  1.630 0.805 2.015 0.895 ;
        RECT  1.835 1.005 1.925 1.325 ;
        RECT  1.830 0.275 1.920 0.535 ;
        RECT  1.460 1.235 1.835 1.325 ;
        RECT  1.155 0.275 1.830 0.375 ;
        RECT  1.345 1.425 1.555 1.545 ;
        RECT  1.505 0.545 1.510 0.715 ;
        RECT  1.415 0.545 1.505 1.145 ;
        RECT  1.285 0.545 1.415 0.650 ;
        RECT  1.350 1.055 1.415 1.145 ;
        RECT  1.260 1.055 1.350 1.335 ;
        RECT  0.450 1.425 1.345 1.525 ;
        RECT  1.065 0.275 1.155 0.660 ;
        RECT  0.780 0.570 1.065 0.660 ;
        RECT  0.685 0.570 0.780 1.155 ;
        RECT  0.670 0.355 0.685 1.155 ;
        RECT  0.575 0.355 0.670 0.660 ;
        RECT  0.540 1.045 0.670 1.155 ;
        RECT  0.450 0.750 0.520 0.920 ;
        RECT  0.360 0.505 0.450 1.525 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.435 0.360 1.525 ;
        RECT  0.075 0.365 0.185 0.595 ;
        RECT  0.075 1.205 0.185 1.525 ;
    END
END DFCSND4

MACRO DFCSNQD1
    CLASS CORE ;
    FOREIGN DFCSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0755 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.890 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.020 0.295 5.150 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0533 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.760 1.290 0.945 ;
        RECT  1.150 0.800 1.180 0.945 ;
        RECT  1.050 0.800 1.150 1.300 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0737 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.710 4.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.180 -0.165 5.200 0.165 ;
        RECT  4.010 -0.165 4.180 0.620 ;
        RECT  2.220 -0.165 4.010 0.165 ;
        RECT  2.050 -0.165 2.220 0.355 ;
        RECT  0.945 -0.165 2.050 0.165 ;
        RECT  0.835 -0.165 0.945 0.480 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.650 1.635 5.200 1.965 ;
        RECT  3.485 1.435 3.650 1.965 ;
        RECT  3.480 1.435 3.485 1.525 ;
        RECT  2.760 1.635 3.485 1.965 ;
        RECT  2.570 1.425 2.760 1.965 ;
        RECT  0.000 1.635 2.570 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.800 0.515 4.910 1.500 ;
        RECT  4.630 0.515 4.800 0.640 ;
        RECT  4.090 1.390 4.800 1.500 ;
        RECT  4.500 0.265 4.630 0.640 ;
        RECT  4.460 0.750 4.570 1.295 ;
        RECT  3.870 1.205 4.460 1.295 ;
        RECT  4.000 1.390 4.090 1.545 ;
        RECT  3.830 1.435 4.000 1.545 ;
        RECT  3.625 1.025 3.955 1.115 ;
        RECT  3.780 1.205 3.870 1.335 ;
        RECT  3.175 1.245 3.780 1.335 ;
        RECT  3.360 0.510 3.695 0.620 ;
        RECT  3.360 1.025 3.625 1.155 ;
        RECT  3.270 0.510 3.360 1.155 ;
        RECT  2.435 0.315 3.350 0.415 ;
        RECT  3.055 0.570 3.270 0.695 ;
        RECT  3.070 0.825 3.175 1.335 ;
        RECT  2.945 0.825 3.070 0.915 ;
        RECT  2.885 1.245 2.975 1.525 ;
        RECT  2.835 0.525 2.945 0.915 ;
        RECT  2.680 1.055 2.940 1.155 ;
        RECT  2.415 1.245 2.885 1.335 ;
        RECT  2.560 0.505 2.680 1.155 ;
        RECT  2.105 1.055 2.560 1.155 ;
        RECT  2.345 0.315 2.435 0.535 ;
        RECT  2.325 1.245 2.415 1.525 ;
        RECT  1.920 0.445 2.345 0.535 ;
        RECT  1.555 1.425 2.325 1.525 ;
        RECT  2.200 0.625 2.315 0.940 ;
        RECT  1.510 0.625 2.200 0.715 ;
        RECT  2.015 0.805 2.105 1.155 ;
        RECT  1.630 0.805 2.015 0.895 ;
        RECT  1.835 1.005 1.925 1.325 ;
        RECT  1.830 0.275 1.920 0.535 ;
        RECT  1.460 1.235 1.835 1.325 ;
        RECT  1.155 0.275 1.830 0.375 ;
        RECT  1.345 1.425 1.555 1.545 ;
        RECT  1.505 0.545 1.510 0.715 ;
        RECT  1.415 0.545 1.505 1.145 ;
        RECT  1.285 0.545 1.415 0.650 ;
        RECT  1.350 1.055 1.415 1.145 ;
        RECT  1.260 1.055 1.350 1.335 ;
        RECT  0.450 1.425 1.345 1.525 ;
        RECT  1.065 0.275 1.155 0.660 ;
        RECT  0.800 0.570 1.065 0.660 ;
        RECT  0.685 0.570 0.800 1.315 ;
        RECT  0.660 0.355 0.685 1.315 ;
        RECT  0.575 0.355 0.660 0.660 ;
        RECT  0.540 1.205 0.660 1.315 ;
        RECT  0.450 0.750 0.520 0.920 ;
        RECT  0.360 0.505 0.450 1.525 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.435 0.360 1.525 ;
        RECT  0.075 0.365 0.185 0.595 ;
        RECT  0.075 1.205 0.185 1.525 ;
    END
END DFCSNQD1

MACRO DFCSNQD2
    CLASS CORE ;
    FOREIGN DFCSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0755 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.890 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.280 5.550 1.495 ;
        RECT  5.355 0.280 5.450 0.660 ;
        RECT  5.350 1.025 5.450 1.495 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0533 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.760 1.290 0.945 ;
        RECT  1.150 0.800 1.180 0.945 ;
        RECT  1.050 0.800 1.150 1.300 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1289 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.920 0.600 5.030 0.910 ;
        RECT  4.550 0.600 4.920 0.690 ;
        RECT  4.420 0.600 4.550 1.100 ;
        RECT  4.100 0.780 4.420 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.190 -0.165 5.800 0.165 ;
        RECT  4.055 -0.165 4.190 0.635 ;
        RECT  2.220 -0.165 4.055 0.165 ;
        RECT  2.050 -0.165 2.220 0.355 ;
        RECT  0.945 -0.165 2.050 0.165 ;
        RECT  0.835 -0.165 0.945 0.480 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.650 1.635 5.800 1.965 ;
        RECT  3.485 1.435 3.650 1.965 ;
        RECT  3.480 1.435 3.485 1.525 ;
        RECT  2.760 1.635 3.485 1.965 ;
        RECT  2.570 1.425 2.760 1.965 ;
        RECT  0.000 1.635 2.570 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.225 0.750 5.300 0.920 ;
        RECT  5.120 0.400 5.225 1.500 ;
        RECT  4.540 0.400 5.120 0.510 ;
        RECT  4.090 1.390 5.120 1.500 ;
        RECT  4.640 0.815 4.810 1.295 ;
        RECT  3.870 1.205 4.640 1.295 ;
        RECT  4.000 1.390 4.090 1.545 ;
        RECT  3.830 1.435 4.000 1.545 ;
        RECT  3.625 1.025 3.955 1.115 ;
        RECT  3.780 1.205 3.870 1.335 ;
        RECT  3.175 1.245 3.780 1.335 ;
        RECT  3.360 0.510 3.700 0.620 ;
        RECT  3.360 1.025 3.625 1.155 ;
        RECT  3.270 0.510 3.360 1.155 ;
        RECT  2.435 0.315 3.350 0.415 ;
        RECT  3.055 0.570 3.270 0.695 ;
        RECT  3.070 0.825 3.175 1.335 ;
        RECT  2.945 0.825 3.070 0.915 ;
        RECT  2.885 1.245 2.975 1.525 ;
        RECT  2.835 0.525 2.945 0.915 ;
        RECT  2.680 1.055 2.940 1.155 ;
        RECT  2.415 1.245 2.885 1.335 ;
        RECT  2.560 0.505 2.680 1.155 ;
        RECT  2.105 1.055 2.560 1.155 ;
        RECT  2.345 0.315 2.435 0.535 ;
        RECT  2.325 1.245 2.415 1.525 ;
        RECT  1.920 0.445 2.345 0.535 ;
        RECT  1.555 1.425 2.325 1.525 ;
        RECT  2.200 0.625 2.315 0.940 ;
        RECT  1.510 0.625 2.200 0.715 ;
        RECT  2.015 0.805 2.105 1.155 ;
        RECT  1.630 0.805 2.015 0.895 ;
        RECT  1.835 1.005 1.925 1.325 ;
        RECT  1.830 0.275 1.920 0.535 ;
        RECT  1.460 1.235 1.835 1.325 ;
        RECT  1.155 0.275 1.830 0.375 ;
        RECT  1.345 1.425 1.555 1.545 ;
        RECT  1.505 0.545 1.510 0.715 ;
        RECT  1.415 0.545 1.505 1.145 ;
        RECT  1.285 0.545 1.415 0.650 ;
        RECT  1.350 1.055 1.415 1.145 ;
        RECT  1.260 1.055 1.350 1.335 ;
        RECT  0.450 1.425 1.345 1.525 ;
        RECT  1.065 0.275 1.155 0.660 ;
        RECT  0.800 0.570 1.065 0.660 ;
        RECT  0.685 0.570 0.800 1.315 ;
        RECT  0.660 0.355 0.685 1.315 ;
        RECT  0.575 0.355 0.660 0.660 ;
        RECT  0.540 1.205 0.660 1.315 ;
        RECT  0.450 0.750 0.520 0.920 ;
        RECT  0.360 0.505 0.450 1.525 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.435 0.360 1.525 ;
        RECT  0.075 0.365 0.185 0.595 ;
        RECT  0.075 1.205 0.185 1.525 ;
    END
END DFCSNQD2

MACRO DFCSNQD4
    CLASS CORE ;
    FOREIGN DFCSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0755 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.890 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.475 6.070 0.660 ;
        RECT  5.850 1.080 6.070 1.300 ;
        RECT  5.530 0.475 5.850 1.300 ;
        RECT  5.365 0.475 5.530 0.660 ;
        RECT  5.345 1.080 5.530 1.300 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0533 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.760 1.290 0.945 ;
        RECT  1.150 0.800 1.180 0.945 ;
        RECT  1.050 0.800 1.150 1.300 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1289 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.945 0.610 5.055 0.910 ;
        RECT  4.550 0.610 4.945 0.700 ;
        RECT  4.430 0.610 4.550 1.100 ;
        RECT  4.100 0.780 4.430 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.225 -0.165 6.400 0.165 ;
        RECT  4.050 -0.165 4.225 0.665 ;
        RECT  2.220 -0.165 4.050 0.165 ;
        RECT  2.050 -0.165 2.220 0.355 ;
        RECT  0.945 -0.165 2.050 0.165 ;
        RECT  0.835 -0.165 0.945 0.480 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.290 1.635 6.400 1.965 ;
        RECT  6.175 1.010 6.290 1.965 ;
        RECT  5.795 1.635 6.175 1.965 ;
        RECT  5.625 1.410 5.795 1.965 ;
        RECT  3.650 1.635 5.625 1.965 ;
        RECT  3.485 1.435 3.650 1.965 ;
        RECT  3.480 1.435 3.485 1.525 ;
        RECT  2.760 1.635 3.485 1.965 ;
        RECT  2.570 1.425 2.760 1.965 ;
        RECT  0.000 1.635 2.570 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.950 0.475 6.070 0.660 ;
        RECT  5.950 1.080 6.070 1.300 ;
        RECT  5.365 0.475 5.450 0.660 ;
        RECT  5.345 1.080 5.450 1.300 ;
        RECT  5.245 0.750 5.330 0.920 ;
        RECT  5.145 0.390 5.245 1.500 ;
        RECT  4.550 0.390 5.145 0.505 ;
        RECT  4.090 1.390 5.145 1.500 ;
        RECT  4.640 0.815 4.810 1.295 ;
        RECT  3.870 1.205 4.640 1.295 ;
        RECT  4.000 1.390 4.090 1.545 ;
        RECT  3.830 1.435 4.000 1.545 ;
        RECT  3.625 1.025 3.955 1.115 ;
        RECT  3.780 1.205 3.870 1.335 ;
        RECT  3.175 1.245 3.780 1.335 ;
        RECT  3.360 0.510 3.695 0.620 ;
        RECT  3.360 1.025 3.625 1.155 ;
        RECT  3.270 0.510 3.360 1.155 ;
        RECT  2.435 0.315 3.350 0.415 ;
        RECT  3.055 0.570 3.270 0.695 ;
        RECT  3.070 0.825 3.175 1.335 ;
        RECT  2.945 0.825 3.070 0.915 ;
        RECT  2.885 1.245 2.975 1.525 ;
        RECT  2.835 0.525 2.945 0.915 ;
        RECT  2.680 1.055 2.940 1.155 ;
        RECT  2.415 1.245 2.885 1.335 ;
        RECT  2.560 0.505 2.680 1.155 ;
        RECT  2.105 1.055 2.560 1.155 ;
        RECT  2.345 0.315 2.435 0.535 ;
        RECT  2.325 1.245 2.415 1.525 ;
        RECT  1.920 0.445 2.345 0.535 ;
        RECT  1.555 1.425 2.325 1.525 ;
        RECT  2.200 0.625 2.315 0.940 ;
        RECT  1.510 0.625 2.200 0.715 ;
        RECT  2.015 0.805 2.105 1.155 ;
        RECT  1.630 0.805 2.015 0.895 ;
        RECT  1.835 1.005 1.925 1.325 ;
        RECT  1.830 0.275 1.920 0.535 ;
        RECT  1.460 1.235 1.835 1.325 ;
        RECT  1.155 0.275 1.830 0.375 ;
        RECT  1.345 1.425 1.555 1.545 ;
        RECT  1.505 0.545 1.510 0.715 ;
        RECT  1.415 0.545 1.505 1.145 ;
        RECT  1.285 0.545 1.415 0.650 ;
        RECT  1.350 1.055 1.415 1.145 ;
        RECT  1.260 1.055 1.350 1.335 ;
        RECT  0.450 1.425 1.345 1.525 ;
        RECT  1.065 0.275 1.155 0.660 ;
        RECT  0.800 0.570 1.065 0.660 ;
        RECT  0.685 0.570 0.800 1.315 ;
        RECT  0.660 0.275 0.685 1.315 ;
        RECT  0.575 0.275 0.660 0.660 ;
        RECT  0.540 1.205 0.660 1.315 ;
        RECT  0.450 0.750 0.520 0.920 ;
        RECT  0.360 0.505 0.450 1.525 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.435 0.360 1.525 ;
        RECT  0.075 0.365 0.185 0.595 ;
        RECT  0.075 1.205 0.185 1.525 ;
    END
END DFCSNQD4

MACRO DFD1
    CLASS CORE ;
    FOREIGN DFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.840 0.285 3.950 1.490 ;
        RECT  3.825 0.285 3.840 0.675 ;
        RECT  3.825 1.050 3.840 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.480 3.555 1.490 ;
        RECT  3.325 0.480 3.450 0.650 ;
        RECT  3.325 0.995 3.450 1.185 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.245 0.920 ;
        RECT  1.050 0.730 1.155 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.670 0.155 1.110 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.885 -0.165 4.000 0.165 ;
        RECT  0.715 -0.165 0.885 0.370 ;
        RECT  0.000 -0.165 0.715 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.735 0.775 3.750 0.945 ;
        RECT  3.645 0.280 3.735 0.945 ;
        RECT  2.850 0.280 3.645 0.370 ;
        RECT  3.235 0.760 3.340 0.890 ;
        RECT  3.145 0.480 3.235 1.525 ;
        RECT  3.070 0.480 3.145 0.660 ;
        RECT  3.120 1.315 3.145 1.525 ;
        RECT  2.625 1.435 3.120 1.525 ;
        RECT  3.030 0.750 3.055 0.930 ;
        RECT  2.940 0.750 3.030 1.345 ;
        RECT  2.420 1.255 2.940 1.345 ;
        RECT  2.760 0.280 2.850 1.165 ;
        RECT  2.575 0.345 2.760 0.520 ;
        RECT  2.560 1.055 2.760 1.165 ;
        RECT  2.485 0.855 2.630 0.965 ;
        RECT  2.395 0.275 2.485 0.965 ;
        RECT  2.305 1.095 2.420 1.345 ;
        RECT  2.235 0.275 2.395 0.365 ;
        RECT  2.075 1.455 2.315 1.545 ;
        RECT  2.300 0.455 2.305 1.345 ;
        RECT  2.195 0.455 2.300 1.185 ;
        RECT  2.065 0.255 2.235 0.365 ;
        RECT  1.995 0.475 2.105 1.315 ;
        RECT  1.995 1.425 2.075 1.545 ;
        RECT  1.105 0.275 2.065 0.365 ;
        RECT  1.700 0.475 1.995 0.600 ;
        RECT  0.410 1.425 1.995 1.525 ;
        RECT  1.815 0.730 1.905 1.315 ;
        RECT  1.485 1.205 1.815 1.315 ;
        RECT  1.585 0.475 1.700 0.940 ;
        RECT  1.375 0.495 1.485 1.315 ;
        RECT  1.200 0.495 1.375 0.585 ;
        RECT  1.190 1.205 1.375 1.315 ;
        RECT  1.005 0.275 1.105 0.580 ;
        RECT  0.795 0.470 1.005 0.580 ;
        RECT  0.685 0.470 0.795 1.190 ;
        RECT  0.535 0.470 0.685 0.640 ;
        RECT  0.525 1.065 0.685 1.190 ;
        RECT  0.410 0.770 0.530 0.940 ;
        RECT  0.310 0.460 0.410 1.525 ;
        RECT  0.180 0.460 0.310 0.560 ;
        RECT  0.075 1.350 0.310 1.525 ;
        RECT  0.080 0.370 0.180 0.560 ;
    END
END DFD1

MACRO DFD2
    CLASS CORE ;
    FOREIGN DFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.280 4.350 1.490 ;
        RECT  4.165 0.280 4.250 0.660 ;
        RECT  4.165 1.040 4.250 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.715 0.495 3.815 1.490 ;
        RECT  3.610 0.495 3.715 0.630 ;
        RECT  3.650 1.040 3.715 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.245 0.920 ;
        RECT  1.050 0.730 1.155 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.670 0.155 1.110 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.885 -0.165 4.600 0.165 ;
        RECT  0.715 -0.165 0.885 0.370 ;
        RECT  0.000 -0.165 0.715 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.015 0.750 4.140 0.920 ;
        RECT  3.925 0.275 4.015 0.920 ;
        RECT  2.740 0.275 3.925 0.385 ;
        RECT  3.445 0.730 3.600 0.920 ;
        RECT  3.335 0.495 3.445 1.475 ;
        RECT  2.940 0.495 3.335 0.605 ;
        RECT  3.165 1.305 3.335 1.475 ;
        RECT  3.090 0.750 3.210 1.205 ;
        RECT  2.940 1.080 3.090 1.205 ;
        RECT  2.830 0.495 2.940 0.940 ;
        RECT  2.850 1.080 2.940 1.525 ;
        RECT  2.515 1.435 2.850 1.525 ;
        RECT  2.650 0.275 2.740 1.335 ;
        RECT  2.585 0.275 2.650 0.675 ;
        RECT  2.630 1.120 2.650 1.335 ;
        RECT  2.485 0.855 2.560 1.025 ;
        RECT  2.425 1.255 2.515 1.525 ;
        RECT  2.395 0.275 2.485 1.025 ;
        RECT  2.420 1.255 2.425 1.345 ;
        RECT  2.305 1.120 2.420 1.345 ;
        RECT  2.235 0.275 2.395 0.365 ;
        RECT  2.075 1.455 2.315 1.545 ;
        RECT  2.300 0.455 2.305 1.345 ;
        RECT  2.195 0.455 2.300 1.210 ;
        RECT  2.065 0.255 2.235 0.365 ;
        RECT  1.995 0.475 2.105 1.315 ;
        RECT  1.995 1.425 2.075 1.545 ;
        RECT  1.105 0.275 2.065 0.365 ;
        RECT  1.700 0.475 1.995 0.600 ;
        RECT  0.410 1.425 1.995 1.525 ;
        RECT  1.815 0.730 1.905 1.315 ;
        RECT  1.485 1.205 1.815 1.315 ;
        RECT  1.585 0.475 1.700 0.940 ;
        RECT  1.375 0.495 1.485 1.315 ;
        RECT  1.200 0.495 1.375 0.585 ;
        RECT  1.190 1.205 1.375 1.315 ;
        RECT  1.005 0.275 1.105 0.580 ;
        RECT  0.795 0.470 1.005 0.580 ;
        RECT  0.685 0.470 0.795 1.190 ;
        RECT  0.535 0.470 0.685 0.640 ;
        RECT  0.525 1.065 0.685 1.190 ;
        RECT  0.410 0.770 0.530 0.940 ;
        RECT  0.310 0.460 0.410 1.525 ;
        RECT  0.180 0.460 0.310 0.560 ;
        RECT  0.075 1.350 0.310 1.525 ;
        RECT  0.080 0.370 0.180 0.560 ;
    END
END DFD2

MACRO DFD4
    CLASS CORE ;
    FOREIGN DFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.495 4.225 0.670 ;
        RECT  4.050 1.040 4.225 1.255 ;
        RECT  3.760 0.495 4.050 1.255 ;
        RECT  3.505 0.495 3.760 0.670 ;
        RECT  3.505 1.040 3.760 1.255 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.310 5.710 0.690 ;
        RECT  5.450 1.110 5.710 1.490 ;
        RECT  5.150 0.310 5.450 1.490 ;
        RECT  5.050 0.310 5.150 0.690 ;
        RECT  5.030 1.110 5.150 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.165 0.710 1.255 0.920 ;
        RECT  1.050 0.710 1.165 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.670 0.155 1.110 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.165 6.000 0.165 ;
        RECT  0.760 -0.165 0.930 0.395 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 6.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.550 0.310 5.710 0.690 ;
        RECT  5.550 1.110 5.710 1.490 ;
        RECT  4.150 0.495 4.225 0.670 ;
        RECT  4.150 1.040 4.225 1.255 ;
        RECT  3.505 0.495 3.660 0.670 ;
        RECT  3.505 1.040 3.660 1.255 ;
        RECT  4.870 0.780 5.060 0.890 ;
        RECT  4.770 0.555 4.870 1.140 ;
        RECT  4.675 0.555 4.770 0.655 ;
        RECT  4.675 1.040 4.770 1.140 ;
        RECT  4.565 0.275 4.675 0.655 ;
        RECT  4.565 1.040 4.675 1.470 ;
        RECT  4.430 0.780 4.660 0.890 ;
        RECT  3.155 0.275 4.565 0.385 ;
        RECT  4.330 0.780 4.430 1.475 ;
        RECT  2.470 1.365 4.330 1.475 ;
        RECT  3.365 0.780 3.625 0.890 ;
        RECT  3.240 0.505 3.365 1.275 ;
        RECT  2.595 0.505 3.240 0.675 ;
        RECT  2.560 1.155 3.240 1.275 ;
        RECT  2.985 0.255 3.155 0.385 ;
        RECT  2.495 0.855 2.570 1.025 ;
        RECT  2.405 0.275 2.495 1.025 ;
        RECT  2.430 1.255 2.470 1.475 ;
        RECT  2.380 1.120 2.430 1.475 ;
        RECT  2.245 0.275 2.405 0.365 ;
        RECT  2.315 1.120 2.380 1.345 ;
        RECT  2.310 0.455 2.315 1.345 ;
        RECT  2.205 0.455 2.310 1.210 ;
        RECT  2.085 1.455 2.270 1.545 ;
        RECT  2.075 0.255 2.245 0.365 ;
        RECT  2.005 0.475 2.115 1.315 ;
        RECT  2.005 1.425 2.085 1.545 ;
        RECT  1.110 0.275 2.075 0.365 ;
        RECT  1.710 0.475 2.005 0.600 ;
        RECT  0.420 1.425 2.005 1.525 ;
        RECT  1.825 0.730 1.915 1.315 ;
        RECT  1.495 1.205 1.825 1.315 ;
        RECT  1.595 0.475 1.710 0.940 ;
        RECT  1.385 0.475 1.495 1.315 ;
        RECT  1.210 0.475 1.385 0.585 ;
        RECT  1.200 1.205 1.385 1.315 ;
        RECT  1.020 0.275 1.110 0.620 ;
        RECT  0.800 0.500 1.020 0.620 ;
        RECT  0.680 0.500 0.800 1.160 ;
        RECT  0.540 0.500 0.680 0.660 ;
        RECT  0.525 1.040 0.680 1.160 ;
        RECT  0.420 0.770 0.570 0.900 ;
        RECT  0.320 0.460 0.420 1.525 ;
        RECT  0.180 0.460 0.320 0.560 ;
        RECT  0.075 1.230 0.320 1.400 ;
        RECT  0.080 0.370 0.180 0.560 ;
    END
END DFD4

MACRO DFKCND1
    CLASS CORE ;
    FOREIGN DFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.275 4.550 1.490 ;
        RECT  4.415 0.275 4.450 0.675 ;
        RECT  4.415 1.045 4.450 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1710 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.555 0.465 3.750 0.575 ;
        RECT  3.555 1.160 3.735 1.290 ;
        RECT  3.445 0.465 3.555 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.770 1.350 0.910 ;
        RECT  1.045 0.495 1.155 0.910 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.180 1.120 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.500 0.955 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.635 4.600 1.965 ;
        RECT  2.130 1.310 2.240 1.965 ;
        RECT  0.000 1.635 2.130 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.310 0.765 4.355 0.955 ;
        RECT  4.215 0.275 4.310 0.955 ;
        RECT  3.190 0.275 4.215 0.365 ;
        RECT  3.905 0.475 4.015 1.265 ;
        RECT  2.845 1.415 3.920 1.525 ;
        RECT  3.665 0.760 3.905 0.910 ;
        RECT  3.080 0.275 3.190 1.305 ;
        RECT  2.875 0.275 2.970 1.275 ;
        RECT  1.990 0.275 2.875 0.365 ;
        RECT  2.845 1.050 2.875 1.275 ;
        RECT  2.755 1.385 2.845 1.525 ;
        RECT  2.755 0.465 2.785 0.800 ;
        RECT  2.665 0.465 2.755 1.525 ;
        RECT  2.635 1.385 2.665 1.525 ;
        RECT  2.480 0.475 2.575 1.220 ;
        RECT  2.375 0.475 2.480 0.605 ;
        RECT  2.110 1.110 2.480 1.220 ;
        RECT  2.270 0.700 2.390 1.005 ;
        RECT  1.890 0.700 2.270 0.790 ;
        RECT  2.000 0.905 2.110 1.220 ;
        RECT  1.580 0.275 1.990 0.385 ;
        RECT  1.850 0.495 1.890 0.790 ;
        RECT  0.425 1.435 1.870 1.525 ;
        RECT  1.740 0.495 1.850 1.270 ;
        RECT  1.675 0.495 1.740 0.625 ;
        RECT  1.590 1.160 1.740 1.270 ;
        RECT  1.470 0.275 1.580 1.060 ;
        RECT  0.775 1.220 1.475 1.330 ;
        RECT  0.745 0.275 1.470 0.385 ;
        RECT  0.685 0.275 0.745 1.130 ;
        RECT  0.655 0.275 0.685 1.330 ;
        RECT  0.550 0.275 0.655 0.485 ;
        RECT  0.575 1.020 0.655 1.330 ;
        RECT  0.425 0.770 0.560 0.900 ;
        RECT  0.335 0.450 0.425 1.525 ;
        RECT  0.185 0.450 0.335 0.560 ;
        RECT  0.290 1.230 0.335 1.525 ;
        RECT  0.075 1.230 0.290 1.410 ;
        RECT  0.075 0.290 0.185 0.560 ;
    END
END DFKCND1

MACRO DFKCND2
    CLASS CORE ;
    FOREIGN DFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.470 3.750 1.295 ;
        RECT  3.515 0.470 3.650 0.580 ;
        RECT  3.515 1.205 3.650 1.295 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.275 4.750 1.490 ;
        RECT  4.565 0.275 4.650 0.675 ;
        RECT  4.565 1.040 4.650 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.770 1.350 0.910 ;
        RECT  1.045 0.495 1.155 0.910 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.180 1.120 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.500 0.955 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.635 5.000 1.965 ;
        RECT  2.130 1.310 2.240 1.965 ;
        RECT  0.000 1.635 2.130 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.780 4.560 0.890 ;
        RECT  4.315 0.575 4.425 1.140 ;
        RECT  4.175 0.575 4.315 0.675 ;
        RECT  4.175 1.040 4.315 1.140 ;
        RECT  3.960 0.780 4.225 0.890 ;
        RECT  4.065 0.275 4.175 0.675 ;
        RECT  4.065 1.040 4.175 1.470 ;
        RECT  3.330 0.275 4.065 0.365 ;
        RECT  3.860 0.780 3.960 1.495 ;
        RECT  2.755 1.385 3.860 1.495 ;
        RECT  3.450 0.730 3.560 1.115 ;
        RECT  3.175 1.025 3.450 1.115 ;
        RECT  3.240 0.275 3.330 0.915 ;
        RECT  3.150 1.025 3.175 1.265 ;
        RECT  3.060 0.290 3.150 1.265 ;
        RECT  2.875 0.275 2.970 1.275 ;
        RECT  1.990 0.275 2.875 0.365 ;
        RECT  2.845 1.050 2.875 1.275 ;
        RECT  2.755 0.465 2.785 0.800 ;
        RECT  2.665 0.465 2.755 1.495 ;
        RECT  2.635 1.385 2.665 1.495 ;
        RECT  2.480 0.475 2.575 1.220 ;
        RECT  2.375 0.475 2.480 0.605 ;
        RECT  2.110 1.110 2.480 1.220 ;
        RECT  2.270 0.700 2.390 1.005 ;
        RECT  1.890 0.700 2.270 0.790 ;
        RECT  2.000 0.905 2.110 1.220 ;
        RECT  1.580 0.275 1.990 0.385 ;
        RECT  1.850 0.495 1.890 0.790 ;
        RECT  0.425 1.435 1.870 1.525 ;
        RECT  1.740 0.495 1.850 1.270 ;
        RECT  1.675 0.495 1.740 0.625 ;
        RECT  1.590 1.160 1.740 1.270 ;
        RECT  1.470 0.275 1.580 1.060 ;
        RECT  0.775 1.220 1.475 1.330 ;
        RECT  0.745 0.275 1.470 0.385 ;
        RECT  0.685 0.275 0.745 1.130 ;
        RECT  0.655 0.275 0.685 1.330 ;
        RECT  0.550 0.275 0.655 0.485 ;
        RECT  0.575 1.020 0.655 1.330 ;
        RECT  0.425 0.770 0.560 0.900 ;
        RECT  0.335 0.450 0.425 1.525 ;
        RECT  0.185 0.450 0.335 0.560 ;
        RECT  0.290 1.230 0.335 1.525 ;
        RECT  0.075 1.230 0.290 1.410 ;
        RECT  0.075 0.290 0.185 0.560 ;
    END
END DFKCND2

MACRO DFKCND4
    CLASS CORE ;
    FOREIGN DFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.470 4.730 0.580 ;
        RECT  4.450 1.155 4.730 1.265 ;
        RECT  4.150 0.470 4.450 1.265 ;
        RECT  4.020 0.470 4.150 0.580 ;
        RECT  4.020 1.155 4.150 1.265 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.120 0.275 6.230 0.675 ;
        RECT  6.120 1.040 6.230 1.470 ;
        RECT  6.050 0.575 6.120 0.675 ;
        RECT  6.050 1.040 6.120 1.140 ;
        RECT  5.750 0.575 6.050 1.140 ;
        RECT  5.710 0.575 5.750 0.675 ;
        RECT  5.710 1.040 5.750 1.140 ;
        RECT  5.600 0.275 5.710 0.675 ;
        RECT  5.600 1.040 5.710 1.470 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.765 1.350 0.910 ;
        RECT  1.045 0.495 1.155 0.910 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.180 1.120 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.500 0.955 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.490 -0.165 6.600 0.165 ;
        RECT  6.380 -0.165 6.490 0.695 ;
        RECT  5.970 -0.165 6.380 0.165 ;
        RECT  5.860 -0.165 5.970 0.475 ;
        RECT  5.450 -0.165 5.860 0.165 ;
        RECT  5.340 -0.165 5.450 0.475 ;
        RECT  0.000 -0.165 5.340 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.490 1.635 6.600 1.965 ;
        RECT  6.380 1.040 6.490 1.965 ;
        RECT  5.970 1.635 6.380 1.965 ;
        RECT  5.860 1.260 5.970 1.965 ;
        RECT  5.450 1.635 5.860 1.965 ;
        RECT  5.340 1.260 5.450 1.965 ;
        RECT  2.250 1.635 5.340 1.965 ;
        RECT  2.140 1.310 2.250 1.965 ;
        RECT  0.000 1.635 2.140 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.150 0.275 6.230 0.675 ;
        RECT  6.150 1.040 6.230 1.470 ;
        RECT  5.600 0.275 5.650 0.675 ;
        RECT  5.600 1.040 5.650 1.470 ;
        RECT  4.550 0.470 4.730 0.580 ;
        RECT  4.550 1.155 4.730 1.265 ;
        RECT  4.020 0.470 4.050 0.580 ;
        RECT  4.020 1.155 4.050 1.265 ;
        RECT  5.460 0.780 5.595 0.890 ;
        RECT  5.350 0.575 5.460 1.140 ;
        RECT  5.190 0.575 5.350 0.675 ;
        RECT  5.190 1.040 5.350 1.140 ;
        RECT  4.925 0.780 5.240 0.890 ;
        RECT  5.080 0.275 5.190 0.675 ;
        RECT  5.080 1.040 5.190 1.470 ;
        RECT  3.430 0.275 5.080 0.365 ;
        RECT  4.825 0.780 4.925 1.495 ;
        RECT  2.785 1.385 4.825 1.495 ;
        RECT  3.660 0.780 3.960 0.890 ;
        RECT  3.660 1.155 3.755 1.265 ;
        RECT  3.550 0.470 3.660 1.265 ;
        RECT  3.150 1.155 3.550 1.265 ;
        RECT  3.320 0.275 3.430 0.935 ;
        RECT  3.060 0.295 3.150 1.265 ;
        RECT  2.875 0.275 2.970 1.265 ;
        RECT  2.395 0.275 2.875 0.365 ;
        RECT  2.675 0.465 2.785 1.495 ;
        RECT  2.645 1.385 2.675 1.495 ;
        RECT  2.495 0.495 2.585 1.220 ;
        RECT  2.375 0.495 2.495 0.605 ;
        RECT  2.135 1.110 2.495 1.220 ;
        RECT  2.305 0.275 2.395 0.405 ;
        RECT  2.270 0.700 2.380 1.005 ;
        RECT  1.580 0.295 2.305 0.405 ;
        RECT  1.900 0.700 2.270 0.790 ;
        RECT  2.020 0.920 2.135 1.220 ;
        RECT  0.425 1.435 1.910 1.525 ;
        RECT  1.790 0.500 1.900 1.270 ;
        RECT  1.675 0.500 1.790 0.635 ;
        RECT  1.590 1.160 1.790 1.270 ;
        RECT  1.470 0.295 1.580 1.060 ;
        RECT  0.775 1.220 1.475 1.330 ;
        RECT  0.745 0.295 1.470 0.405 ;
        RECT  0.655 0.295 0.745 1.130 ;
        RECT  0.535 0.545 0.655 0.655 ;
        RECT  0.535 1.020 0.655 1.130 ;
        RECT  0.425 0.770 0.560 0.900 ;
        RECT  0.335 0.450 0.425 1.525 ;
        RECT  0.185 0.450 0.335 0.560 ;
        RECT  0.185 1.435 0.335 1.525 ;
        RECT  0.075 0.290 0.185 0.560 ;
        RECT  0.075 1.270 0.185 1.525 ;
    END
END DFKCND4

MACRO DFKCNQD1
    CLASS CORE ;
    FOREIGN DFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.275 3.950 1.490 ;
        RECT  3.825 0.275 3.850 0.660 ;
        RECT  3.815 1.020 3.850 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0443 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.220 0.710 1.350 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.160 1.110 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0445 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.750 1.020 0.920 ;
        RECT  0.850 0.660 0.950 1.090 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.215 -0.165 4.000 0.165 ;
        RECT  3.080 -0.165 3.215 0.355 ;
        RECT  0.985 -0.165 3.080 0.165 ;
        RECT  0.815 -0.165 0.985 0.355 ;
        RECT  0.000 -0.165 0.815 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.205 1.635 4.000 1.965 ;
        RECT  2.030 1.355 2.205 1.965 ;
        RECT  0.000 1.635 2.030 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.670 0.750 3.760 0.920 ;
        RECT  3.570 0.485 3.670 1.420 ;
        RECT  3.070 0.485 3.570 0.615 ;
        RECT  3.260 1.310 3.570 1.420 ;
        RECT  3.290 0.745 3.420 1.160 ;
        RECT  3.125 1.070 3.290 1.160 ;
        RECT  3.035 1.070 3.125 1.495 ;
        RECT  2.980 0.485 3.070 0.960 ;
        RECT  2.665 1.395 3.035 1.495 ;
        RECT  2.845 0.275 2.880 0.950 ;
        RECT  2.790 0.275 2.845 1.285 ;
        RECT  2.575 0.275 2.790 0.365 ;
        RECT  2.755 0.835 2.790 1.285 ;
        RECT  2.665 0.465 2.700 0.660 ;
        RECT  2.575 0.465 2.665 1.495 ;
        RECT  2.365 0.255 2.575 0.365 ;
        RECT  2.545 1.395 2.575 1.495 ;
        RECT  2.380 0.475 2.485 1.245 ;
        RECT  2.235 0.475 2.380 0.585 ;
        RECT  2.040 1.135 2.380 1.245 ;
        RECT  1.860 0.275 2.365 0.365 ;
        RECT  2.175 0.700 2.280 1.005 ;
        RECT  1.740 0.700 2.175 0.790 ;
        RECT  1.920 0.880 2.040 1.245 ;
        RECT  1.645 0.255 1.860 0.365 ;
        RECT  1.610 1.420 1.835 1.545 ;
        RECT  1.695 0.465 1.740 0.790 ;
        RECT  1.565 0.465 1.695 1.330 ;
        RECT  1.275 0.275 1.645 0.365 ;
        RECT  0.465 1.420 1.610 1.525 ;
        RECT  0.785 1.190 1.455 1.300 ;
        RECT  1.185 0.275 1.275 0.535 ;
        RECT  0.690 0.445 1.185 0.535 ;
        RECT  0.600 0.285 0.690 1.215 ;
        RECT  0.585 0.285 0.600 0.530 ;
        RECT  0.585 1.045 0.600 1.215 ;
        RECT  0.465 0.750 0.510 0.920 ;
        RECT  0.375 0.510 0.465 1.525 ;
        RECT  0.195 0.510 0.375 0.600 ;
        RECT  0.075 1.220 0.375 1.390 ;
        RECT  0.070 0.285 0.195 0.600 ;
    END
END DFKCNQD1

MACRO DFKCNQD2
    CLASS CORE ;
    FOREIGN DFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 0.510 4.150 1.120 ;
        RECT  4.075 0.275 4.080 1.120 ;
        RECT  4.050 0.275 4.075 1.490 ;
        RECT  3.955 0.275 4.050 0.675 ;
        RECT  3.945 1.020 4.050 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0443 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.220 0.710 1.350 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.160 1.110 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0445 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.750 1.020 0.920 ;
        RECT  0.850 0.660 0.950 1.090 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.335 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.335 0.445 ;
        RECT  3.810 -0.165 4.215 0.165 ;
        RECT  3.680 -0.165 3.810 0.465 ;
        RECT  3.240 -0.165 3.680 0.165 ;
        RECT  3.110 -0.165 3.240 0.465 ;
        RECT  0.985 -0.165 3.110 0.165 ;
        RECT  0.815 -0.165 0.985 0.355 ;
        RECT  0.000 -0.165 0.815 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.335 1.635 4.400 1.965 ;
        RECT  4.215 1.260 4.335 1.965 ;
        RECT  3.810 1.635 4.215 1.965 ;
        RECT  3.680 1.335 3.810 1.965 ;
        RECT  3.260 1.635 3.680 1.965 ;
        RECT  3.130 1.335 3.260 1.965 ;
        RECT  2.205 1.635 3.130 1.965 ;
        RECT  2.030 1.355 2.205 1.965 ;
        RECT  0.000 1.635 2.030 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.810 0.780 3.950 0.890 ;
        RECT  3.700 0.575 3.810 1.140 ;
        RECT  3.535 0.575 3.700 0.670 ;
        RECT  3.535 1.040 3.700 1.140 ;
        RECT  3.270 0.780 3.585 0.890 ;
        RECT  3.425 0.275 3.535 0.670 ;
        RECT  3.425 1.040 3.535 1.470 ;
        RECT  3.080 0.575 3.425 0.670 ;
        RECT  3.170 0.780 3.270 1.180 ;
        RECT  3.040 1.090 3.170 1.180 ;
        RECT  2.970 0.575 3.080 0.960 ;
        RECT  2.950 1.090 3.040 1.495 ;
        RECT  2.665 1.395 2.950 1.495 ;
        RECT  2.845 0.275 2.880 0.950 ;
        RECT  2.790 0.275 2.845 1.285 ;
        RECT  2.575 0.275 2.790 0.365 ;
        RECT  2.755 0.835 2.790 1.285 ;
        RECT  2.665 0.465 2.700 0.660 ;
        RECT  2.575 0.465 2.665 1.495 ;
        RECT  2.365 0.255 2.575 0.365 ;
        RECT  2.545 1.395 2.575 1.495 ;
        RECT  2.380 0.475 2.485 1.245 ;
        RECT  2.235 0.475 2.380 0.585 ;
        RECT  2.040 1.135 2.380 1.245 ;
        RECT  1.860 0.275 2.365 0.365 ;
        RECT  2.175 0.700 2.280 1.005 ;
        RECT  1.740 0.700 2.175 0.790 ;
        RECT  1.920 0.880 2.040 1.245 ;
        RECT  1.645 0.255 1.860 0.365 ;
        RECT  1.610 1.420 1.835 1.545 ;
        RECT  1.695 0.465 1.740 0.790 ;
        RECT  1.565 0.465 1.695 1.330 ;
        RECT  1.275 0.275 1.645 0.365 ;
        RECT  0.465 1.420 1.610 1.525 ;
        RECT  0.785 1.190 1.455 1.300 ;
        RECT  1.185 0.275 1.275 0.535 ;
        RECT  0.690 0.445 1.185 0.535 ;
        RECT  0.600 0.285 0.690 1.215 ;
        RECT  0.585 0.285 0.600 0.530 ;
        RECT  0.585 1.045 0.600 1.215 ;
        RECT  0.465 0.750 0.510 0.920 ;
        RECT  0.375 0.510 0.465 1.525 ;
        RECT  0.195 0.510 0.375 0.600 ;
        RECT  0.075 1.220 0.375 1.390 ;
        RECT  0.070 0.285 0.195 0.600 ;
    END
END DFKCNQD2

MACRO DFKCNQD4
    CLASS CORE ;
    FOREIGN DFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.310 4.495 0.675 ;
        RECT  4.250 1.060 4.475 1.430 ;
        RECT  3.950 0.310 4.250 1.430 ;
        RECT  3.825 0.310 3.950 0.675 ;
        RECT  3.850 1.060 3.950 1.430 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0443 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.360 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.160 1.110 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0445 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.750 1.030 0.920 ;
        RECT  0.850 0.660 0.960 1.090 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.725 -0.165 4.800 0.165 ;
        RECT  4.615 -0.165 4.725 0.685 ;
        RECT  3.220 -0.165 4.615 0.165 ;
        RECT  3.080 -0.165 3.220 0.465 ;
        RECT  0.995 -0.165 3.080 0.165 ;
        RECT  0.825 -0.165 0.995 0.355 ;
        RECT  0.000 -0.165 0.825 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.725 1.635 4.800 1.965 ;
        RECT  4.615 1.050 4.725 1.965 ;
        RECT  2.215 1.635 4.615 1.965 ;
        RECT  2.040 1.355 2.215 1.965 ;
        RECT  0.000 1.635 2.040 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.350 0.310 4.495 0.675 ;
        RECT  4.350 1.060 4.475 1.430 ;
        RECT  3.710 0.765 3.840 0.920 ;
        RECT  3.605 0.575 3.710 1.140 ;
        RECT  3.465 0.575 3.605 0.670 ;
        RECT  3.465 1.040 3.605 1.140 ;
        RECT  3.265 0.780 3.495 0.890 ;
        RECT  3.355 0.275 3.465 0.670 ;
        RECT  3.355 1.040 3.465 1.470 ;
        RECT  3.080 0.575 3.355 0.670 ;
        RECT  3.170 0.780 3.265 1.495 ;
        RECT  2.675 1.395 3.170 1.495 ;
        RECT  2.980 0.575 3.080 0.960 ;
        RECT  2.800 0.275 2.890 1.285 ;
        RECT  2.585 0.275 2.800 0.365 ;
        RECT  2.765 1.060 2.800 1.285 ;
        RECT  2.675 0.465 2.710 0.660 ;
        RECT  2.585 0.465 2.675 1.495 ;
        RECT  2.375 0.255 2.585 0.365 ;
        RECT  2.555 1.395 2.585 1.495 ;
        RECT  2.390 0.475 2.495 1.245 ;
        RECT  2.245 0.475 2.390 0.585 ;
        RECT  2.050 1.135 2.390 1.245 ;
        RECT  1.870 0.275 2.375 0.365 ;
        RECT  2.185 0.700 2.290 1.005 ;
        RECT  1.750 0.700 2.185 0.790 ;
        RECT  1.930 0.880 2.050 1.245 ;
        RECT  1.655 0.255 1.870 0.365 ;
        RECT  1.620 1.420 1.845 1.545 ;
        RECT  1.705 0.465 1.750 0.790 ;
        RECT  1.575 0.465 1.705 1.330 ;
        RECT  1.285 0.275 1.655 0.365 ;
        RECT  0.465 1.420 1.620 1.525 ;
        RECT  0.795 1.190 1.465 1.300 ;
        RECT  1.195 0.275 1.285 0.535 ;
        RECT  0.690 0.445 1.195 0.535 ;
        RECT  0.600 0.285 0.690 1.215 ;
        RECT  0.585 0.285 0.600 0.660 ;
        RECT  0.585 1.045 0.600 1.215 ;
        RECT  0.465 0.750 0.510 0.920 ;
        RECT  0.375 0.510 0.465 1.525 ;
        RECT  0.195 0.510 0.375 0.600 ;
        RECT  0.075 1.220 0.375 1.390 ;
        RECT  0.070 0.365 0.195 0.600 ;
    END
END DFKCNQD4

MACRO DFKCSND1
    CLASS CORE ;
    FOREIGN DFKCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0310 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.660 0.160 1.090 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.275 5.150 1.490 ;
        RECT  5.020 0.275 5.050 0.675 ;
        RECT  5.005 1.040 5.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.485 4.750 1.100 ;
        RECT  4.525 0.485 4.650 0.655 ;
        RECT  4.635 1.000 4.650 1.100 ;
        RECT  4.515 1.000 4.635 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.995 0.770 1.225 ;
        RECT  0.650 0.995 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.710 1.550 1.090 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0328 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.635 1.260 1.135 ;
        RECT  0.550 0.635 1.170 0.725 ;
        RECT  0.910 1.025 1.170 1.135 ;
        RECT  0.440 0.310 0.550 0.725 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.855 1.635 5.200 1.965 ;
        RECT  2.855 1.210 3.000 1.320 ;
        RECT  2.745 1.210 2.855 1.965 ;
        RECT  0.000 1.635 2.745 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.930 0.750 4.950 0.940 ;
        RECT  4.840 0.275 4.930 0.940 ;
        RECT  3.835 0.275 4.840 0.385 ;
        RECT  4.425 0.765 4.540 0.895 ;
        RECT  4.365 0.510 4.425 1.300 ;
        RECT  4.335 0.510 4.365 1.450 ;
        RECT  4.015 0.510 4.335 0.620 ;
        RECT  4.250 1.210 4.335 1.450 ;
        RECT  4.155 0.730 4.245 1.100 ;
        RECT  4.095 1.010 4.155 1.100 ;
        RECT  4.000 1.010 4.095 1.495 ;
        RECT  3.925 0.510 4.015 0.895 ;
        RECT  3.445 1.395 4.000 1.495 ;
        RECT  3.745 0.275 3.835 1.195 ;
        RECT  3.565 0.275 3.655 1.305 ;
        RECT  3.390 0.275 3.565 0.365 ;
        RECT  3.535 1.135 3.565 1.305 ;
        RECT  3.445 0.465 3.475 0.975 ;
        RECT  3.355 0.465 3.445 1.495 ;
        RECT  3.220 0.265 3.390 0.365 ;
        RECT  3.175 0.495 3.265 1.320 ;
        RECT  3.150 0.275 3.220 0.365 ;
        RECT  2.855 0.495 3.175 0.605 ;
        RECT  3.090 1.210 3.175 1.320 ;
        RECT  3.060 0.275 3.150 0.405 ;
        RECT  2.975 0.795 3.085 1.120 ;
        RECT  2.485 0.295 3.060 0.405 ;
        RECT  2.530 1.030 2.975 1.120 ;
        RECT  2.745 0.495 2.855 0.940 ;
        RECT  2.520 0.500 2.530 1.120 ;
        RECT  2.420 0.500 2.520 1.365 ;
        RECT  2.395 1.140 2.420 1.365 ;
        RECT  2.175 0.545 2.285 1.165 ;
        RECT  0.945 1.400 2.270 1.510 ;
        RECT  2.080 0.265 2.250 0.410 ;
        RECT  1.850 0.545 2.175 0.655 ;
        RECT  1.850 1.055 2.175 1.165 ;
        RECT  1.020 0.310 2.080 0.410 ;
        RECT  1.750 0.770 1.915 0.900 ;
        RECT  1.660 0.500 1.750 1.310 ;
        RECT  1.370 0.500 1.660 0.620 ;
        RECT  1.370 1.200 1.660 1.310 ;
        RECT  0.910 0.815 1.080 0.925 ;
        RECT  0.850 0.310 1.020 0.545 ;
        RECT  0.840 1.335 0.945 1.510 ;
        RECT  0.530 0.815 0.910 0.905 ;
        RECT  0.395 0.815 0.530 1.345 ;
        RECT  0.340 0.815 0.395 0.925 ;
        RECT  0.185 1.255 0.395 1.345 ;
        RECT  0.250 0.335 0.340 0.925 ;
        RECT  0.045 0.335 0.250 0.435 ;
        RECT  0.075 1.255 0.185 1.515 ;
    END
END DFKCSND1

MACRO DFKCSND2
    CLASS CORE ;
    FOREIGN DFKCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.750 0.180 0.920 ;
        RECT  0.050 0.660 0.150 1.090 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.575 5.150 1.215 ;
        RECT  4.975 0.575 5.050 0.675 ;
        RECT  4.815 1.105 5.050 1.215 ;
        RECT  4.865 0.275 4.975 0.675 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.365 0.275 5.550 0.690 ;
        RECT  5.350 1.105 5.505 1.215 ;
        RECT  5.350 0.575 5.365 0.690 ;
        RECT  5.250 0.575 5.350 1.215 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0247 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.035 0.860 1.225 ;
        RECT  0.650 1.035 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.570 1.090 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0297 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.635 1.350 1.195 ;
        RECT  0.590 0.635 1.240 0.725 ;
        RECT  0.980 1.085 1.240 1.195 ;
        RECT  0.480 0.535 0.590 0.725 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.470 -0.165 5.800 0.165 ;
        RECT  0.360 -0.165 0.470 0.340 ;
        RECT  0.000 -0.165 0.360 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.930 1.635 5.800 1.965 ;
        RECT  2.930 1.210 3.075 1.320 ;
        RECT  2.820 1.210 2.930 1.965 ;
        RECT  0.475 1.635 2.820 1.965 ;
        RECT  0.365 1.455 0.475 1.965 ;
        RECT  0.000 1.635 0.365 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.595 0.780 5.685 1.475 ;
        RECT  5.460 0.780 5.595 0.890 ;
        RECT  4.585 1.375 5.595 1.475 ;
        RECT  4.775 0.780 4.940 0.890 ;
        RECT  4.675 0.275 4.775 0.890 ;
        RECT  3.940 0.275 4.675 0.385 ;
        RECT  4.495 0.510 4.585 1.475 ;
        RECT  4.130 0.510 4.495 0.620 ;
        RECT  4.315 1.365 4.495 1.475 ;
        RECT  4.295 0.730 4.405 1.255 ;
        RECT  4.170 1.155 4.295 1.255 ;
        RECT  4.080 1.155 4.170 1.495 ;
        RECT  4.030 0.510 4.130 0.935 ;
        RECT  3.550 1.385 4.080 1.495 ;
        RECT  3.940 1.025 3.975 1.265 ;
        RECT  3.850 0.275 3.940 1.265 ;
        RECT  3.670 0.275 3.760 1.265 ;
        RECT  3.225 0.275 3.670 0.365 ;
        RECT  3.640 1.055 3.670 1.265 ;
        RECT  3.550 0.465 3.580 0.655 ;
        RECT  3.460 0.465 3.550 1.495 ;
        RECT  3.430 1.390 3.460 1.495 ;
        RECT  3.280 0.495 3.370 1.320 ;
        RECT  2.955 0.495 3.280 0.605 ;
        RECT  3.165 1.210 3.280 1.320 ;
        RECT  3.135 0.275 3.225 0.405 ;
        RECT  3.090 0.795 3.190 1.120 ;
        RECT  2.575 0.295 3.135 0.405 ;
        RECT  2.605 1.030 3.090 1.120 ;
        RECT  2.840 0.495 2.955 0.940 ;
        RECT  2.595 0.500 2.605 1.120 ;
        RECT  2.495 0.500 2.595 1.365 ;
        RECT  2.470 1.140 2.495 1.365 ;
        RECT  2.140 0.830 2.405 0.940 ;
        RECT  1.270 0.310 2.370 0.415 ;
        RECT  1.330 1.400 2.345 1.510 ;
        RECT  2.050 0.590 2.140 1.195 ;
        RECT  1.930 0.590 2.050 0.700 ;
        RECT  1.930 1.085 2.050 1.195 ;
        RECT  1.820 0.840 1.955 0.970 ;
        RECT  1.730 0.505 1.820 1.310 ;
        RECT  1.440 0.505 1.730 0.600 ;
        RECT  1.440 1.200 1.730 1.310 ;
        RECT  1.220 1.335 1.330 1.510 ;
        RECT  1.180 0.310 1.270 0.545 ;
        RECT  0.865 1.335 1.220 1.445 ;
        RECT  0.900 0.445 1.180 0.545 ;
        RECT  0.550 0.835 1.150 0.925 ;
        RECT  0.440 0.835 0.550 1.345 ;
        RECT  0.370 0.835 0.440 0.925 ;
        RECT  0.185 1.255 0.440 1.345 ;
        RECT  0.280 0.450 0.370 0.925 ;
        RECT  0.045 0.450 0.280 0.550 ;
        RECT  0.075 1.255 0.185 1.515 ;
    END
END DFKCSND2

MACRO DFKCSND4
    CLASS CORE ;
    FOREIGN DFKCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0310 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.660 0.160 1.090 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.400 5.880 0.600 ;
        RECT  5.650 1.055 5.880 1.255 ;
        RECT  5.350 0.400 5.650 1.255 ;
        RECT  5.220 0.400 5.350 0.600 ;
        RECT  5.170 1.055 5.350 1.255 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 1.060 6.880 1.450 ;
        RECT  6.650 0.370 6.850 0.615 ;
        RECT  6.350 0.370 6.650 1.450 ;
        RECT  6.170 0.370 6.350 0.615 ;
        RECT  6.200 1.060 6.350 1.450 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.995 0.770 1.225 ;
        RECT  0.650 0.995 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.710 1.550 1.090 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0328 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.635 1.260 1.135 ;
        RECT  0.550 0.635 1.170 0.725 ;
        RECT  0.910 1.025 1.170 1.135 ;
        RECT  0.440 0.310 0.550 0.725 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.120 -0.165 7.200 0.165 ;
        RECT  6.990 -0.165 7.120 0.695 ;
        RECT  0.000 -0.165 6.990 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.120 1.635 7.200 1.965 ;
        RECT  6.990 1.040 7.120 1.965 ;
        RECT  2.830 1.635 6.990 1.965 ;
        RECT  2.830 1.210 2.975 1.320 ;
        RECT  2.720 1.210 2.830 1.965 ;
        RECT  0.000 1.635 2.720 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.750 1.060 6.880 1.450 ;
        RECT  6.750 0.370 6.850 0.615 ;
        RECT  6.170 0.370 6.250 0.615 ;
        RECT  6.200 1.060 6.250 1.450 ;
        RECT  5.790 0.400 5.880 0.600 ;
        RECT  5.790 1.055 5.880 1.255 ;
        RECT  5.220 0.400 5.310 0.600 ;
        RECT  5.170 1.055 5.310 1.255 ;
        RECT  6.080 0.780 6.260 0.890 ;
        RECT  5.970 0.780 6.080 1.465 ;
        RECT  4.940 1.365 5.970 1.465 ;
        RECT  5.130 0.780 5.260 0.890 ;
        RECT  5.030 0.275 5.130 0.890 ;
        RECT  4.345 0.275 5.030 0.385 ;
        RECT  4.850 0.510 4.940 1.465 ;
        RECT  4.550 0.510 4.850 0.620 ;
        RECT  4.670 1.355 4.850 1.465 ;
        RECT  4.650 0.730 4.760 1.125 ;
        RECT  4.545 1.025 4.650 1.125 ;
        RECT  4.440 0.510 4.550 0.890 ;
        RECT  4.445 1.025 4.545 1.495 ;
        RECT  3.450 1.385 4.445 1.495 ;
        RECT  3.945 0.780 4.440 0.890 ;
        RECT  4.235 1.025 4.350 1.275 ;
        RECT  4.235 0.275 4.345 0.675 ;
        RECT  3.835 0.275 4.235 0.380 ;
        RECT  3.835 1.185 4.235 1.275 ;
        RECT  3.740 0.275 3.835 1.275 ;
        RECT  3.540 0.275 3.650 1.295 ;
        RECT  3.365 0.275 3.540 0.365 ;
        RECT  3.340 0.465 3.450 1.495 ;
        RECT  3.195 0.265 3.365 0.365 ;
        RECT  3.150 0.495 3.240 1.320 ;
        RECT  3.125 0.275 3.195 0.365 ;
        RECT  2.830 0.495 3.150 0.605 ;
        RECT  3.065 1.210 3.150 1.320 ;
        RECT  3.035 0.275 3.125 0.405 ;
        RECT  2.950 0.795 3.060 1.120 ;
        RECT  2.460 0.295 3.035 0.405 ;
        RECT  2.505 1.030 2.950 1.120 ;
        RECT  2.720 0.495 2.830 0.940 ;
        RECT  2.495 0.500 2.505 1.120 ;
        RECT  2.395 0.500 2.495 1.365 ;
        RECT  2.370 1.140 2.395 1.365 ;
        RECT  1.020 0.310 2.270 0.410 ;
        RECT  2.150 0.545 2.260 1.165 ;
        RECT  0.945 1.400 2.245 1.510 ;
        RECT  1.835 0.545 2.150 0.655 ;
        RECT  1.835 1.055 2.150 1.165 ;
        RECT  1.735 0.770 1.900 0.900 ;
        RECT  1.645 0.500 1.735 1.310 ;
        RECT  1.355 0.500 1.645 0.620 ;
        RECT  1.355 1.200 1.645 1.310 ;
        RECT  0.910 0.815 1.080 0.925 ;
        RECT  0.850 0.310 1.020 0.545 ;
        RECT  0.840 1.335 0.945 1.510 ;
        RECT  0.530 0.815 0.910 0.905 ;
        RECT  0.395 0.815 0.530 1.345 ;
        RECT  0.340 0.815 0.395 0.925 ;
        RECT  0.185 1.255 0.395 1.345 ;
        RECT  0.250 0.335 0.340 0.925 ;
        RECT  0.045 0.335 0.250 0.435 ;
        RECT  0.075 1.255 0.185 1.515 ;
    END
END DFKCSND4

MACRO DFKSND1
    CLASS CORE ;
    FOREIGN DFKSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.710 1.030 0.920 ;
        RECT  0.850 0.710 0.950 1.090 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.575 4.550 1.100 ;
        RECT  4.425 0.575 4.450 0.675 ;
        RECT  4.425 1.000 4.450 1.100 ;
        RECT  4.315 0.475 4.425 0.675 ;
        RECT  4.315 1.000 4.425 1.265 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.275 4.950 1.490 ;
        RECT  4.815 0.275 4.850 0.675 ;
        RECT  4.820 1.040 4.850 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0377 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.700 1.550 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.750 0.280 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.625 1.635 5.000 1.965 ;
        RECT  2.625 1.215 2.745 1.315 ;
        RECT  2.515 1.215 2.625 1.965 ;
        RECT  0.000 1.635 2.515 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.730 0.750 4.760 0.940 ;
        RECT  4.640 0.750 4.730 1.475 ;
        RECT  4.220 1.375 4.640 1.475 ;
        RECT  3.600 0.275 4.330 0.385 ;
        RECT  4.130 0.510 4.220 1.475 ;
        RECT  3.790 0.510 4.130 0.620 ;
        RECT  3.975 1.365 4.130 1.475 ;
        RECT  3.930 0.730 4.040 1.255 ;
        RECT  3.865 1.155 3.930 1.255 ;
        RECT  3.775 1.155 3.865 1.495 ;
        RECT  3.690 0.510 3.790 0.935 ;
        RECT  3.215 1.385 3.775 1.495 ;
        RECT  3.600 1.025 3.635 1.275 ;
        RECT  3.510 0.275 3.600 1.275 ;
        RECT  3.305 0.275 3.400 1.265 ;
        RECT  0.700 0.275 3.305 0.375 ;
        RECT  3.105 0.465 3.215 1.495 ;
        RECT  3.075 1.385 3.105 1.495 ;
        RECT  2.925 0.495 3.015 1.300 ;
        RECT  2.565 0.495 2.925 0.605 ;
        RECT  2.835 1.190 2.925 1.300 ;
        RECT  2.700 0.795 2.810 1.100 ;
        RECT  2.340 1.010 2.700 1.100 ;
        RECT  2.450 0.495 2.565 0.920 ;
        RECT  1.910 1.405 2.405 1.515 ;
        RECT  2.250 0.510 2.340 1.315 ;
        RECT  2.065 0.510 2.250 0.620 ;
        RECT  2.020 1.205 2.250 1.315 ;
        RECT  1.910 0.730 2.010 0.840 ;
        RECT  1.730 0.500 1.955 0.610 ;
        RECT  1.820 0.730 1.910 1.515 ;
        RECT  0.470 1.425 1.820 1.515 ;
        RECT  1.640 0.500 1.730 1.315 ;
        RECT  1.300 0.500 1.640 0.610 ;
        RECT  1.495 1.205 1.640 1.315 ;
        RECT  1.210 0.750 1.285 0.920 ;
        RECT  1.120 0.500 1.210 1.315 ;
        RECT  0.805 0.500 1.120 0.600 ;
        RECT  0.800 1.200 1.120 1.315 ;
        RECT  0.610 0.275 0.700 1.280 ;
        RECT  0.580 0.275 0.610 0.585 ;
        RECT  0.575 1.070 0.610 1.280 ;
        RECT  0.470 0.750 0.520 0.920 ;
        RECT  0.370 0.475 0.470 1.515 ;
        RECT  0.185 0.475 0.370 0.585 ;
        RECT  0.185 1.425 0.370 1.515 ;
        RECT  0.075 0.375 0.185 0.585 ;
        RECT  0.075 1.210 0.185 1.515 ;
    END
END DFKSND1

MACRO DFKSND2
    CLASS CORE ;
    FOREIGN DFKSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.710 1.030 0.920 ;
        RECT  0.850 0.710 0.950 1.090 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.575 4.750 1.215 ;
        RECT  4.575 0.575 4.650 0.675 ;
        RECT  4.415 1.105 4.650 1.215 ;
        RECT  4.465 0.275 4.575 0.675 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.965 0.275 5.150 0.690 ;
        RECT  4.950 1.105 5.105 1.215 ;
        RECT  4.950 0.575 4.965 0.690 ;
        RECT  4.850 0.575 4.950 1.215 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0377 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.700 1.550 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.750 0.280 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.545 1.635 5.400 1.965 ;
        RECT  2.545 1.225 2.685 1.335 ;
        RECT  2.445 1.225 2.545 1.965 ;
        RECT  0.000 1.635 2.445 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.195 0.780 5.285 1.475 ;
        RECT  5.060 0.780 5.195 0.890 ;
        RECT  4.185 1.375 5.195 1.475 ;
        RECT  4.375 0.780 4.540 0.890 ;
        RECT  4.275 0.275 4.375 0.890 ;
        RECT  3.540 0.275 4.275 0.385 ;
        RECT  4.095 0.510 4.185 1.475 ;
        RECT  3.730 0.510 4.095 0.620 ;
        RECT  3.915 1.365 4.095 1.475 ;
        RECT  3.895 0.730 4.005 1.255 ;
        RECT  3.825 1.155 3.895 1.255 ;
        RECT  3.735 1.155 3.825 1.495 ;
        RECT  3.150 1.385 3.735 1.495 ;
        RECT  3.630 0.510 3.730 0.895 ;
        RECT  3.540 0.985 3.575 1.175 ;
        RECT  3.450 0.275 3.540 1.175 ;
        RECT  3.270 0.275 3.360 1.295 ;
        RECT  0.700 0.275 3.270 0.365 ;
        RECT  3.240 1.085 3.270 1.295 ;
        RECT  3.150 0.465 3.180 0.655 ;
        RECT  3.060 0.465 3.150 1.495 ;
        RECT  2.880 0.495 2.970 1.325 ;
        RECT  2.545 0.495 2.880 0.605 ;
        RECT  2.795 1.215 2.880 1.325 ;
        RECT  2.690 0.795 2.790 1.125 ;
        RECT  2.305 1.035 2.690 1.125 ;
        RECT  2.435 0.495 2.545 0.945 ;
        RECT  1.920 1.415 2.320 1.515 ;
        RECT  2.215 0.480 2.305 1.125 ;
        RECT  2.065 0.480 2.215 0.590 ;
        RECT  2.120 1.035 2.215 1.125 ;
        RECT  2.010 1.035 2.120 1.320 ;
        RECT  1.730 0.455 1.955 0.550 ;
        RECT  1.820 0.660 1.920 1.515 ;
        RECT  0.470 1.425 1.820 1.515 ;
        RECT  1.640 0.455 1.730 1.315 ;
        RECT  1.300 0.485 1.640 0.595 ;
        RECT  1.495 1.205 1.640 1.315 ;
        RECT  1.210 0.780 1.330 0.890 ;
        RECT  1.120 0.500 1.210 1.315 ;
        RECT  0.805 0.500 1.120 0.600 ;
        RECT  0.800 1.200 1.120 1.315 ;
        RECT  0.610 0.275 0.700 1.280 ;
        RECT  0.580 0.275 0.610 0.585 ;
        RECT  0.575 1.070 0.610 1.280 ;
        RECT  0.470 0.750 0.520 0.920 ;
        RECT  0.370 0.475 0.470 1.515 ;
        RECT  0.185 0.475 0.370 0.585 ;
        RECT  0.185 1.425 0.370 1.515 ;
        RECT  0.075 0.375 0.185 0.585 ;
        RECT  0.075 1.210 0.185 1.515 ;
    END
END DFKSND2

MACRO DFKSND4
    CLASS CORE ;
    FOREIGN DFKSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.710 1.030 0.920 ;
        RECT  0.850 0.710 0.950 1.090 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 1.090 5.640 1.200 ;
        RECT  5.480 0.275 5.590 0.675 ;
        RECT  5.450 0.575 5.480 0.675 ;
        RECT  5.150 0.575 5.450 1.200 ;
        RECT  5.070 0.575 5.150 0.675 ;
        RECT  4.910 1.090 5.150 1.200 ;
        RECT  4.960 0.275 5.070 0.675 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.520 0.275 6.630 0.675 ;
        RECT  6.520 1.050 6.630 1.470 ;
        RECT  6.450 0.575 6.520 0.675 ;
        RECT  6.450 1.050 6.520 1.160 ;
        RECT  6.150 0.575 6.450 1.160 ;
        RECT  6.110 0.575 6.150 0.675 ;
        RECT  6.110 1.050 6.150 1.160 ;
        RECT  6.000 0.275 6.110 0.675 ;
        RECT  6.000 1.050 6.110 1.470 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0377 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.700 1.550 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.750 0.280 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.890 -0.165 7.000 0.165 ;
        RECT  6.780 -0.165 6.890 0.685 ;
        RECT  6.370 -0.165 6.780 0.165 ;
        RECT  6.260 -0.165 6.370 0.465 ;
        RECT  5.850 -0.165 6.260 0.165 ;
        RECT  5.740 -0.165 5.850 0.465 ;
        RECT  5.330 -0.165 5.740 0.165 ;
        RECT  5.220 -0.165 5.330 0.465 ;
        RECT  0.000 -0.165 5.220 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.890 1.635 7.000 1.965 ;
        RECT  6.780 1.050 6.890 1.965 ;
        RECT  6.370 1.635 6.780 1.965 ;
        RECT  6.260 1.270 6.370 1.965 ;
        RECT  2.545 1.635 6.260 1.965 ;
        RECT  2.545 1.225 2.685 1.335 ;
        RECT  2.445 1.225 2.545 1.965 ;
        RECT  0.000 1.635 2.445 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.550 0.275 6.630 0.675 ;
        RECT  6.550 1.050 6.630 1.470 ;
        RECT  6.000 0.275 6.050 0.675 ;
        RECT  6.000 1.050 6.050 1.470 ;
        RECT  5.550 1.090 5.640 1.200 ;
        RECT  5.550 0.275 5.590 0.675 ;
        RECT  4.960 0.275 5.050 0.675 ;
        RECT  4.910 1.090 5.050 1.200 ;
        RECT  5.840 0.780 6.050 0.890 ;
        RECT  5.750 0.780 5.840 1.410 ;
        RECT  4.660 1.310 5.750 1.410 ;
        RECT  4.870 0.780 5.035 0.890 ;
        RECT  4.770 0.275 4.870 0.890 ;
        RECT  4.050 0.275 4.770 0.385 ;
        RECT  4.570 0.510 4.660 1.410 ;
        RECT  4.270 0.510 4.570 0.620 ;
        RECT  4.390 1.300 4.570 1.410 ;
        RECT  4.370 0.730 4.480 1.190 ;
        RECT  4.300 1.090 4.370 1.190 ;
        RECT  4.210 1.090 4.300 1.495 ;
        RECT  4.160 0.510 4.270 0.890 ;
        RECT  3.150 1.385 4.210 1.495 ;
        RECT  3.655 0.780 4.160 0.890 ;
        RECT  3.965 0.985 4.075 1.250 ;
        RECT  3.940 0.275 4.050 0.675 ;
        RECT  3.575 0.985 3.965 1.095 ;
        RECT  3.550 0.565 3.940 0.675 ;
        RECT  3.540 0.985 3.575 1.175 ;
        RECT  3.540 0.445 3.550 0.675 ;
        RECT  3.450 0.445 3.540 1.175 ;
        RECT  3.270 0.275 3.360 1.295 ;
        RECT  0.700 0.275 3.270 0.365 ;
        RECT  3.240 1.085 3.270 1.295 ;
        RECT  3.150 0.465 3.180 0.655 ;
        RECT  3.060 0.465 3.150 1.495 ;
        RECT  2.880 0.495 2.970 1.325 ;
        RECT  2.545 0.495 2.880 0.605 ;
        RECT  2.795 1.215 2.880 1.325 ;
        RECT  2.690 0.795 2.790 1.125 ;
        RECT  2.305 1.035 2.690 1.125 ;
        RECT  2.435 0.495 2.545 0.945 ;
        RECT  1.920 1.415 2.320 1.515 ;
        RECT  2.215 0.480 2.305 1.125 ;
        RECT  2.065 0.480 2.215 0.590 ;
        RECT  2.120 1.035 2.215 1.125 ;
        RECT  2.010 1.035 2.120 1.320 ;
        RECT  1.730 0.455 1.955 0.550 ;
        RECT  1.820 0.660 1.920 1.515 ;
        RECT  0.470 1.425 1.820 1.515 ;
        RECT  1.640 0.455 1.730 1.315 ;
        RECT  1.300 0.485 1.640 0.595 ;
        RECT  1.495 1.205 1.640 1.315 ;
        RECT  1.210 0.780 1.330 0.890 ;
        RECT  1.120 0.500 1.210 1.315 ;
        RECT  0.805 0.500 1.120 0.600 ;
        RECT  0.800 1.200 1.120 1.315 ;
        RECT  0.610 0.275 0.700 1.280 ;
        RECT  0.580 0.275 0.610 0.540 ;
        RECT  0.575 1.070 0.610 1.280 ;
        RECT  0.470 0.750 0.520 0.920 ;
        RECT  0.370 0.475 0.470 1.515 ;
        RECT  0.185 0.475 0.370 0.585 ;
        RECT  0.185 1.425 0.370 1.515 ;
        RECT  0.075 0.375 0.185 0.585 ;
        RECT  0.075 1.210 0.185 1.515 ;
    END
END DFKSND4

MACRO DFNCND1
    CLASS CORE ;
    FOREIGN DFNCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.285 4.755 1.490 ;
        RECT  4.625 0.285 4.650 0.675 ;
        RECT  4.625 1.040 4.650 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1430 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.305 4.355 1.125 ;
        RECT  4.065 0.305 4.245 0.415 ;
        RECT  4.075 1.030 4.245 1.125 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0366 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.270 0.910 ;
        RECT  1.050 0.730 1.155 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.750 0.200 0.940 ;
        RECT  0.045 0.650 0.155 1.110 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0651 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.490 3.755 0.890 ;
        RECT  3.445 0.710 3.650 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 -0.165 4.800 0.165 ;
        RECT  3.390 -0.165 3.560 0.600 ;
        RECT  2.045 -0.165 3.390 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.930 -0.165 1.915 0.165 ;
        RECT  0.760 -0.165 0.930 0.415 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.635 4.800 1.965 ;
        RECT  0.820 1.395 0.940 1.505 ;
        RECT  0.720 1.395 0.820 1.965 ;
        RECT  0.000 1.635 0.720 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.535 0.775 4.560 0.945 ;
        RECT  4.445 0.775 4.535 1.315 ;
        RECT  3.160 1.225 4.445 1.315 ;
        RECT  3.990 0.780 4.135 0.890 ;
        RECT  3.960 0.505 3.990 0.890 ;
        RECT  3.860 0.505 3.960 1.135 ;
        RECT  3.350 1.025 3.860 1.135 ;
        RECT  3.630 1.445 3.855 1.535 ;
        RECT  3.540 1.405 3.630 1.535 ;
        RECT  2.970 1.405 3.540 1.495 ;
        RECT  3.250 0.735 3.350 1.135 ;
        RECT  3.100 0.525 3.300 0.625 ;
        RECT  3.225 0.735 3.250 0.945 ;
        RECT  3.100 1.035 3.160 1.315 ;
        RECT  2.890 0.275 3.120 0.435 ;
        RECT  3.060 0.525 3.100 1.315 ;
        RECT  3.010 0.525 3.060 1.125 ;
        RECT  2.800 0.665 3.010 0.775 ;
        RECT  2.900 1.215 2.970 1.495 ;
        RECT  2.880 0.945 2.900 1.495 ;
        RECT  2.225 0.275 2.890 0.365 ;
        RECT  2.790 0.945 2.880 1.320 ;
        RECT  2.675 0.945 2.790 1.045 ;
        RECT  2.620 1.430 2.790 1.545 ;
        RECT  2.565 0.455 2.675 1.045 ;
        RECT  2.425 1.170 2.670 1.280 ;
        RECT  1.120 1.430 2.620 1.520 ;
        RECT  2.315 0.455 2.425 1.280 ;
        RECT  1.725 1.010 2.315 1.110 ;
        RECT  2.135 0.275 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.770 1.220 2.135 1.340 ;
        RECT  1.460 0.720 2.095 0.820 ;
        RECT  1.470 1.220 1.770 1.315 ;
        RECT  1.615 0.910 1.725 1.110 ;
        RECT  1.570 0.265 1.660 0.605 ;
        RECT  1.335 0.265 1.570 0.375 ;
        RECT  1.380 0.510 1.460 1.110 ;
        RECT  1.360 0.510 1.380 1.320 ;
        RECT  1.215 0.510 1.360 0.620 ;
        RECT  1.290 1.020 1.360 1.320 ;
        RECT  1.210 1.210 1.290 1.320 ;
        RECT  1.030 1.210 1.120 1.520 ;
        RECT  0.790 1.210 1.030 1.305 ;
        RECT  0.680 0.535 0.790 1.305 ;
        RECT  0.525 0.535 0.680 0.645 ;
        RECT  0.525 1.045 0.680 1.155 ;
        RECT  0.410 0.750 0.530 0.920 ;
        RECT  0.310 0.440 0.410 1.330 ;
        RECT  0.185 0.440 0.310 0.540 ;
        RECT  0.185 1.220 0.310 1.330 ;
        RECT  0.075 0.330 0.185 0.540 ;
        RECT  0.075 1.220 0.185 1.455 ;
    END
END DFNCND1

MACRO DFNCND2
    CLASS CORE ;
    FOREIGN DFNCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.150 1.090 5.290 1.220 ;
        RECT  5.150 0.285 5.240 0.675 ;
        RECT  5.050 0.285 5.150 1.220 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.565 4.950 1.220 ;
        RECT  4.750 0.565 4.850 0.690 ;
        RECT  4.580 1.090 4.850 1.220 ;
        RECT  4.630 0.285 4.750 0.690 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0366 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.270 0.910 ;
        RECT  1.050 0.730 1.155 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.750 0.200 0.940 ;
        RECT  0.045 0.650 0.155 1.110 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.1015 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.700 3.750 0.900 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.500 -0.165 5.600 0.165 ;
        RECT  5.390 -0.165 5.500 0.590 ;
        RECT  3.560 -0.165 5.390 0.165 ;
        RECT  3.390 -0.165 3.560 0.590 ;
        RECT  2.045 -0.165 3.390 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.930 -0.165 1.915 0.165 ;
        RECT  0.760 -0.165 0.930 0.415 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.635 5.600 1.965 ;
        RECT  0.820 1.395 0.940 1.505 ;
        RECT  0.720 1.395 0.820 1.965 ;
        RECT  0.000 1.635 0.720 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.380 0.730 5.490 1.430 ;
        RECT  4.105 1.340 5.380 1.430 ;
        RECT  4.400 0.780 4.740 0.890 ;
        RECT  4.300 0.495 4.400 1.135 ;
        RECT  3.850 0.495 4.300 0.605 ;
        RECT  3.350 1.025 4.300 1.135 ;
        RECT  3.985 1.225 4.105 1.430 ;
        RECT  3.160 1.225 3.985 1.315 ;
        RECT  3.630 1.435 3.865 1.545 ;
        RECT  3.540 1.405 3.630 1.545 ;
        RECT  2.970 1.405 3.540 1.495 ;
        RECT  3.250 0.735 3.350 1.135 ;
        RECT  3.100 0.525 3.300 0.625 ;
        RECT  3.225 0.735 3.250 0.945 ;
        RECT  3.100 1.035 3.160 1.315 ;
        RECT  2.890 0.275 3.120 0.435 ;
        RECT  3.060 0.525 3.100 1.315 ;
        RECT  3.010 0.525 3.060 1.125 ;
        RECT  2.800 0.665 3.010 0.775 ;
        RECT  2.900 1.215 2.970 1.495 ;
        RECT  2.880 0.945 2.900 1.495 ;
        RECT  2.225 0.275 2.890 0.365 ;
        RECT  2.790 0.945 2.880 1.320 ;
        RECT  2.675 0.945 2.790 1.045 ;
        RECT  2.620 1.430 2.790 1.545 ;
        RECT  2.565 0.455 2.675 1.045 ;
        RECT  2.425 1.200 2.670 1.310 ;
        RECT  1.120 1.430 2.620 1.520 ;
        RECT  2.315 0.455 2.425 1.310 ;
        RECT  1.725 1.010 2.315 1.110 ;
        RECT  2.135 0.275 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.770 1.220 2.135 1.340 ;
        RECT  1.460 0.720 2.095 0.820 ;
        RECT  1.470 1.220 1.770 1.315 ;
        RECT  1.615 0.910 1.725 1.110 ;
        RECT  1.570 0.265 1.660 0.605 ;
        RECT  1.335 0.265 1.570 0.375 ;
        RECT  1.380 0.510 1.460 1.110 ;
        RECT  1.360 0.510 1.380 1.320 ;
        RECT  1.215 0.510 1.360 0.620 ;
        RECT  1.290 1.020 1.360 1.320 ;
        RECT  1.210 1.210 1.290 1.320 ;
        RECT  1.030 1.210 1.120 1.520 ;
        RECT  0.790 1.210 1.030 1.305 ;
        RECT  0.680 0.535 0.790 1.305 ;
        RECT  0.525 0.535 0.680 0.645 ;
        RECT  0.525 1.045 0.680 1.155 ;
        RECT  0.410 0.750 0.530 0.920 ;
        RECT  0.310 0.440 0.410 1.330 ;
        RECT  0.185 0.440 0.310 0.540 ;
        RECT  0.185 1.220 0.310 1.330 ;
        RECT  0.075 0.330 0.185 0.540 ;
        RECT  0.075 1.220 0.185 1.455 ;
    END
END DFNCND2

MACRO DFNCND4
    CLASS CORE ;
    FOREIGN DFNCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.285 6.750 0.675 ;
        RECT  6.650 1.040 6.750 1.500 ;
        RECT  6.565 0.285 6.650 1.500 ;
        RECT  6.350 0.575 6.565 1.150 ;
        RECT  6.175 0.575 6.350 0.675 ;
        RECT  6.175 1.040 6.350 1.150 ;
        RECT  6.065 0.285 6.175 0.675 ;
        RECT  6.065 1.040 6.175 1.500 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.285 5.750 0.675 ;
        RECT  5.650 1.090 5.720 1.220 ;
        RECT  5.565 0.285 5.650 1.220 ;
        RECT  5.350 0.565 5.565 1.220 ;
        RECT  5.175 0.565 5.350 0.675 ;
        RECT  5.015 1.090 5.350 1.220 ;
        RECT  5.065 0.285 5.175 0.675 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0366 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.730 1.270 0.910 ;
        RECT  1.050 0.730 1.155 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.750 0.200 0.940 ;
        RECT  0.045 0.650 0.155 1.110 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.1013 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.700 4.150 0.900 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.925 -0.165 7.000 0.165 ;
        RECT  4.805 -0.165 4.925 0.675 ;
        RECT  3.930 -0.165 4.805 0.165 ;
        RECT  3.760 -0.165 3.930 0.590 ;
        RECT  3.330 -0.165 3.760 0.165 ;
        RECT  3.200 -0.165 3.330 0.445 ;
        RECT  2.045 -0.165 3.200 0.165 ;
        RECT  1.915 -0.165 2.045 0.405 ;
        RECT  0.935 -0.165 1.915 0.165 ;
        RECT  0.760 -0.165 0.935 0.415 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.635 7.000 1.965 ;
        RECT  0.820 1.395 0.940 1.505 ;
        RECT  0.720 1.395 0.820 1.965 ;
        RECT  0.000 1.635 0.720 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.175 0.575 6.250 0.675 ;
        RECT  6.175 1.040 6.250 1.150 ;
        RECT  6.065 0.285 6.175 0.675 ;
        RECT  6.065 1.040 6.175 1.500 ;
        RECT  5.175 0.565 5.250 0.675 ;
        RECT  5.015 1.090 5.250 1.220 ;
        RECT  5.065 0.285 5.175 0.675 ;
        RECT  5.935 0.780 6.200 0.890 ;
        RECT  5.825 0.780 5.935 1.430 ;
        RECT  4.540 1.340 5.825 1.430 ;
        RECT  4.725 0.780 5.175 0.890 ;
        RECT  4.715 0.780 4.725 1.135 ;
        RECT  4.615 0.495 4.715 1.135 ;
        RECT  4.250 0.495 4.615 0.605 ;
        RECT  3.500 1.025 4.615 1.135 ;
        RECT  4.420 1.225 4.540 1.430 ;
        RECT  3.160 1.225 4.420 1.315 ;
        RECT  4.065 1.435 4.300 1.545 ;
        RECT  3.975 1.405 4.065 1.545 ;
        RECT  2.970 1.405 3.975 1.495 ;
        RECT  3.160 0.535 3.635 0.625 ;
        RECT  3.390 0.735 3.500 1.135 ;
        RECT  3.060 0.535 3.160 1.315 ;
        RECT  2.910 0.275 3.110 0.435 ;
        RECT  2.800 0.665 3.060 0.775 ;
        RECT  2.900 1.215 2.970 1.495 ;
        RECT  2.225 0.275 2.910 0.365 ;
        RECT  2.880 0.945 2.900 1.495 ;
        RECT  2.790 0.945 2.880 1.320 ;
        RECT  2.675 0.945 2.790 1.065 ;
        RECT  2.620 1.430 2.790 1.545 ;
        RECT  2.565 0.455 2.675 1.065 ;
        RECT  2.425 1.200 2.670 1.310 ;
        RECT  1.120 1.430 2.620 1.520 ;
        RECT  2.315 0.455 2.425 1.310 ;
        RECT  1.725 1.010 2.315 1.110 ;
        RECT  2.135 0.275 2.225 0.605 ;
        RECT  2.095 0.720 2.205 0.920 ;
        RECT  1.660 0.515 2.135 0.605 ;
        RECT  1.770 1.220 2.135 1.340 ;
        RECT  1.460 0.720 2.095 0.820 ;
        RECT  1.470 1.220 1.770 1.320 ;
        RECT  1.615 0.910 1.725 1.110 ;
        RECT  1.570 0.265 1.660 0.605 ;
        RECT  1.335 0.265 1.570 0.375 ;
        RECT  1.380 0.510 1.460 1.110 ;
        RECT  1.360 0.510 1.380 1.320 ;
        RECT  1.215 0.510 1.360 0.620 ;
        RECT  1.290 1.020 1.360 1.320 ;
        RECT  1.210 1.210 1.290 1.320 ;
        RECT  1.030 1.210 1.120 1.520 ;
        RECT  0.790 1.210 1.030 1.305 ;
        RECT  0.680 0.535 0.790 1.305 ;
        RECT  0.525 0.535 0.680 0.645 ;
        RECT  0.525 1.045 0.680 1.155 ;
        RECT  0.410 0.750 0.530 0.920 ;
        RECT  0.310 0.440 0.410 1.330 ;
        RECT  0.185 0.440 0.310 0.540 ;
        RECT  0.185 1.220 0.310 1.330 ;
        RECT  0.075 0.330 0.185 0.540 ;
        RECT  0.075 1.220 0.185 1.455 ;
    END
END DFNCND4

MACRO DFNCSND1
    CLASS CORE ;
    FOREIGN DFNCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0793 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.780 4.730 0.900 ;
        RECT  4.450 0.500 4.550 0.900 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.275 5.550 1.490 ;
        RECT  5.420 0.275 5.450 0.675 ;
        RECT  5.420 1.045 5.450 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1430 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.495 5.150 1.320 ;
        RECT  4.865 0.495 5.050 0.605 ;
        RECT  4.865 1.210 5.050 1.320 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0510 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.270 0.945 ;
        RECT  1.050 0.700 1.150 1.090 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.700 4.150 0.900 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.110 -0.165 5.600 0.165 ;
        RECT  1.940 -0.165 2.110 0.355 ;
        RECT  0.000 -0.165 1.940 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.635 5.600 1.965 ;
        RECT  4.180 1.190 4.290 1.965 ;
        RECT  4.050 1.190 4.180 1.300 ;
        RECT  3.695 1.635 4.180 1.965 ;
        RECT  3.500 1.435 3.695 1.965 ;
        RECT  2.745 1.635 3.500 1.965 ;
        RECT  2.575 1.410 2.745 1.965 ;
        RECT  0.955 1.635 2.575 1.965 ;
        RECT  0.785 1.395 0.955 1.965 ;
        RECT  0.000 1.635 0.785 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.330 0.750 5.360 0.920 ;
        RECT  5.240 0.290 5.330 1.520 ;
        RECT  4.765 0.290 5.240 0.380 ;
        RECT  4.745 1.420 5.240 1.520 ;
        RECT  4.850 0.730 4.960 1.100 ;
        RECT  4.340 0.995 4.850 1.100 ;
        RECT  4.655 0.290 4.765 0.630 ;
        RECT  4.645 1.190 4.745 1.520 ;
        RECT  3.505 0.290 4.655 0.380 ;
        RECT  4.385 1.190 4.645 1.300 ;
        RECT  4.240 0.490 4.340 1.100 ;
        RECT  3.610 0.490 4.240 0.600 ;
        RECT  3.940 0.995 4.240 1.100 ;
        RECT  3.830 0.995 3.940 1.205 ;
        RECT  3.610 0.730 3.710 1.345 ;
        RECT  3.185 1.255 3.610 1.345 ;
        RECT  3.415 0.290 3.505 1.125 ;
        RECT  3.025 0.530 3.415 0.655 ;
        RECT  3.315 0.995 3.415 1.125 ;
        RECT  2.305 0.305 3.325 0.415 ;
        RECT  3.095 0.855 3.185 1.345 ;
        RECT  2.915 0.855 3.095 0.945 ;
        RECT  2.880 1.230 2.990 1.525 ;
        RECT  2.660 1.035 2.975 1.140 ;
        RECT  2.790 0.515 2.915 0.945 ;
        RECT  2.200 1.230 2.880 1.320 ;
        RECT  2.530 0.515 2.660 1.140 ;
        RECT  2.125 1.035 2.530 1.140 ;
        RECT  2.215 0.625 2.325 0.905 ;
        RECT  2.215 0.305 2.305 0.535 ;
        RECT  1.815 0.445 2.215 0.535 ;
        RECT  1.455 0.625 2.215 0.715 ;
        RECT  2.110 1.230 2.200 1.525 ;
        RECT  2.035 0.805 2.125 1.140 ;
        RECT  1.150 1.425 2.110 1.525 ;
        RECT  1.560 0.805 2.035 0.895 ;
        RECT  1.815 0.985 1.945 1.335 ;
        RECT  1.725 0.275 1.815 0.535 ;
        RECT  1.545 1.165 1.815 1.335 ;
        RECT  0.450 0.275 1.725 0.375 ;
        RECT  1.450 0.485 1.455 0.715 ;
        RECT  1.360 0.485 1.450 1.305 ;
        RECT  1.205 0.485 1.360 0.595 ;
        RECT  1.240 1.195 1.360 1.305 ;
        RECT  1.050 1.180 1.150 1.525 ;
        RECT  0.800 1.180 1.050 1.275 ;
        RECT  0.690 0.570 0.800 1.275 ;
        RECT  0.685 0.570 0.690 0.660 ;
        RECT  0.540 1.095 0.690 1.275 ;
        RECT  0.575 0.470 0.685 0.660 ;
        RECT  0.450 0.750 0.530 0.920 ;
        RECT  0.360 0.275 0.450 1.380 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.290 0.360 1.380 ;
        RECT  0.075 0.385 0.185 0.595 ;
        RECT  0.075 1.290 0.185 1.500 ;
    END
END DFNCSND1

MACRO DFNCSND2
    CLASS CORE ;
    FOREIGN DFNCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0887 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.900 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.985 0.290 6.150 1.490 ;
        RECT  5.950 0.290 5.985 0.675 ;
        RECT  5.950 1.110 5.985 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 0.490 5.630 1.490 ;
        RECT  5.440 0.490 5.530 0.690 ;
        RECT  5.440 1.065 5.530 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0510 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.270 0.945 ;
        RECT  1.050 0.700 1.150 1.090 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.1063 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 5.150 0.900 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.055 -0.165 6.400 0.165 ;
        RECT  3.945 -0.165 4.055 0.440 ;
        RECT  2.110 -0.165 3.945 0.165 ;
        RECT  1.940 -0.165 2.110 0.355 ;
        RECT  0.000 -0.165 1.940 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.290 1.635 6.400 1.965 ;
        RECT  5.180 1.265 5.290 1.965 ;
        RECT  4.255 1.635 5.180 1.965 ;
        RECT  4.065 1.505 4.255 1.965 ;
        RECT  2.745 1.635 4.065 1.965 ;
        RECT  2.575 1.410 2.745 1.965 ;
        RECT  0.955 1.635 2.575 1.965 ;
        RECT  0.785 1.395 0.955 1.965 ;
        RECT  0.000 1.635 0.785 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.830 0.750 5.875 0.920 ;
        RECT  5.740 0.290 5.830 0.920 ;
        RECT  4.255 0.290 5.740 0.380 ;
        RECT  5.350 0.780 5.440 0.890 ;
        RECT  5.260 0.490 5.350 1.155 ;
        RECT  4.510 0.490 5.260 0.600 ;
        RECT  5.030 1.045 5.260 1.155 ;
        RECT  4.920 1.045 5.030 1.485 ;
        RECT  4.650 0.730 4.760 1.395 ;
        RECT  3.185 1.305 4.650 1.395 ;
        RECT  4.400 0.490 4.510 1.195 ;
        RECT  4.020 0.730 4.400 0.900 ;
        RECT  4.165 0.290 4.255 0.620 ;
        RECT  3.930 0.530 4.165 0.620 ;
        RECT  3.930 1.015 4.020 1.125 ;
        RECT  3.840 0.530 3.930 1.125 ;
        RECT  3.285 0.530 3.840 0.620 ;
        RECT  3.295 1.015 3.840 1.125 ;
        RECT  2.305 0.305 3.325 0.415 ;
        RECT  3.025 0.530 3.285 0.655 ;
        RECT  3.095 0.855 3.185 1.395 ;
        RECT  2.915 0.855 3.095 0.945 ;
        RECT  2.880 1.230 2.990 1.525 ;
        RECT  2.660 1.035 2.975 1.140 ;
        RECT  2.790 0.515 2.915 0.945 ;
        RECT  2.200 1.230 2.880 1.320 ;
        RECT  2.530 0.515 2.660 1.140 ;
        RECT  2.125 1.035 2.530 1.140 ;
        RECT  2.215 0.625 2.325 0.905 ;
        RECT  2.215 0.305 2.305 0.535 ;
        RECT  1.815 0.445 2.215 0.535 ;
        RECT  1.455 0.625 2.215 0.715 ;
        RECT  2.110 1.230 2.200 1.525 ;
        RECT  2.035 0.805 2.125 1.140 ;
        RECT  1.150 1.425 2.110 1.525 ;
        RECT  1.560 0.805 2.035 0.895 ;
        RECT  1.815 0.985 1.945 1.335 ;
        RECT  1.725 0.275 1.815 0.535 ;
        RECT  1.545 1.165 1.815 1.335 ;
        RECT  0.450 0.275 1.725 0.375 ;
        RECT  1.450 0.485 1.455 0.715 ;
        RECT  1.360 0.485 1.450 1.305 ;
        RECT  1.205 0.485 1.360 0.595 ;
        RECT  1.240 1.195 1.360 1.305 ;
        RECT  1.050 1.180 1.150 1.525 ;
        RECT  0.800 1.180 1.050 1.275 ;
        RECT  0.690 0.570 0.800 1.275 ;
        RECT  0.685 0.570 0.690 0.660 ;
        RECT  0.540 1.095 0.690 1.275 ;
        RECT  0.575 0.470 0.685 0.660 ;
        RECT  0.450 0.750 0.530 0.920 ;
        RECT  0.360 0.275 0.450 1.380 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.290 0.360 1.380 ;
        RECT  0.075 0.385 0.185 0.595 ;
        RECT  0.075 1.290 0.185 1.500 ;
    END
END DFNCSND2

MACRO DFNCSND4
    CLASS CORE ;
    FOREIGN DFNCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0887 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.900 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.750 0.305 7.050 1.435 ;
        RECT  6.440 0.305 6.750 0.675 ;
        RECT  6.440 1.045 6.750 1.435 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.490 6.050 0.670 ;
        RECT  5.850 1.065 6.050 1.435 ;
        RECT  5.550 0.490 5.850 1.435 ;
        RECT  5.450 0.490 5.550 0.670 ;
        RECT  5.450 1.065 5.550 1.435 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0510 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.270 0.945 ;
        RECT  1.050 0.700 1.150 1.090 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.705 0.250 0.920 ;
        RECT  0.050 0.705 0.150 1.095 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.1063 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 5.150 0.900 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.310 -0.165 7.400 0.165 ;
        RECT  7.200 -0.165 7.310 0.695 ;
        RECT  4.055 -0.165 7.200 0.165 ;
        RECT  3.945 -0.165 4.055 0.440 ;
        RECT  2.110 -0.165 3.945 0.165 ;
        RECT  1.940 -0.165 2.110 0.355 ;
        RECT  0.000 -0.165 1.940 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.310 1.635 7.400 1.965 ;
        RECT  7.200 1.045 7.310 1.965 ;
        RECT  5.290 1.635 7.200 1.965 ;
        RECT  5.180 1.265 5.290 1.965 ;
        RECT  4.255 1.635 5.180 1.965 ;
        RECT  4.065 1.505 4.255 1.965 ;
        RECT  2.745 1.635 4.065 1.965 ;
        RECT  2.575 1.410 2.745 1.965 ;
        RECT  0.955 1.635 2.575 1.965 ;
        RECT  0.785 1.395 0.955 1.965 ;
        RECT  0.000 1.635 0.785 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.440 0.305 6.650 0.675 ;
        RECT  6.440 1.045 6.650 1.435 ;
        RECT  5.950 0.490 6.050 0.670 ;
        RECT  5.950 1.065 6.050 1.435 ;
        RECT  6.250 0.780 6.600 0.890 ;
        RECT  6.160 0.290 6.250 0.890 ;
        RECT  4.255 0.290 6.160 0.380 ;
        RECT  5.350 0.780 5.440 0.890 ;
        RECT  5.260 0.490 5.350 1.155 ;
        RECT  4.510 0.490 5.260 0.600 ;
        RECT  5.030 1.045 5.260 1.155 ;
        RECT  4.920 1.045 5.030 1.485 ;
        RECT  4.650 0.730 4.760 1.395 ;
        RECT  3.185 1.305 4.650 1.395 ;
        RECT  4.400 0.490 4.510 1.195 ;
        RECT  4.020 0.730 4.400 0.900 ;
        RECT  4.165 0.290 4.255 0.620 ;
        RECT  3.930 0.530 4.165 0.620 ;
        RECT  3.930 1.015 4.020 1.125 ;
        RECT  3.840 0.530 3.930 1.125 ;
        RECT  3.285 0.530 3.840 0.620 ;
        RECT  3.295 1.015 3.840 1.125 ;
        RECT  2.305 0.305 3.325 0.415 ;
        RECT  3.025 0.530 3.285 0.655 ;
        RECT  3.095 0.855 3.185 1.395 ;
        RECT  2.915 0.855 3.095 0.945 ;
        RECT  2.880 1.230 2.990 1.525 ;
        RECT  2.660 1.035 2.975 1.140 ;
        RECT  2.790 0.515 2.915 0.945 ;
        RECT  2.200 1.230 2.880 1.320 ;
        RECT  2.530 0.515 2.660 1.140 ;
        RECT  2.125 1.035 2.530 1.140 ;
        RECT  2.215 0.625 2.325 0.905 ;
        RECT  2.215 0.305 2.305 0.535 ;
        RECT  1.815 0.445 2.215 0.535 ;
        RECT  1.455 0.625 2.215 0.715 ;
        RECT  2.110 1.230 2.200 1.525 ;
        RECT  2.035 0.805 2.125 1.140 ;
        RECT  1.150 1.425 2.110 1.525 ;
        RECT  1.560 0.805 2.035 0.895 ;
        RECT  1.815 0.985 1.945 1.335 ;
        RECT  1.725 0.275 1.815 0.535 ;
        RECT  1.545 1.165 1.815 1.335 ;
        RECT  0.450 0.275 1.725 0.375 ;
        RECT  1.450 0.485 1.455 0.715 ;
        RECT  1.360 0.485 1.450 1.305 ;
        RECT  1.205 0.485 1.360 0.595 ;
        RECT  1.240 1.195 1.360 1.305 ;
        RECT  1.050 1.180 1.150 1.525 ;
        RECT  0.800 1.180 1.050 1.275 ;
        RECT  0.690 0.570 0.800 1.275 ;
        RECT  0.685 0.570 0.690 0.660 ;
        RECT  0.540 1.095 0.690 1.275 ;
        RECT  0.575 0.470 0.685 0.660 ;
        RECT  0.450 0.750 0.530 0.920 ;
        RECT  0.360 0.275 0.450 1.380 ;
        RECT  0.185 0.505 0.360 0.595 ;
        RECT  0.185 1.290 0.360 1.380 ;
        RECT  0.075 0.385 0.185 0.595 ;
        RECT  0.075 1.290 0.185 1.500 ;
    END
END DFNCSND4

MACRO DFND1
    CLASS CORE ;
    FOREIGN DFND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.275 4.150 1.490 ;
        RECT  4.020 0.275 4.050 0.675 ;
        RECT  4.015 1.040 4.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.485 3.750 1.150 ;
        RECT  3.515 0.485 3.650 0.675 ;
        RECT  3.625 1.040 3.650 1.150 ;
        RECT  3.515 1.040 3.625 1.480 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.700 1.300 0.900 ;
        RECT  1.050 0.500 1.150 0.900 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 4.200 0.165 ;
        RECT  0.835 -0.165 0.945 0.670 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 1.635 4.200 1.965 ;
        RECT  0.835 1.305 0.945 1.965 ;
        RECT  0.000 1.635 0.835 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.930 0.750 3.960 0.920 ;
        RECT  3.840 0.275 3.930 0.920 ;
        RECT  2.790 0.275 3.840 0.375 ;
        RECT  3.425 0.780 3.540 0.890 ;
        RECT  3.365 0.525 3.425 1.150 ;
        RECT  3.335 0.525 3.365 1.480 ;
        RECT  2.975 0.525 3.335 0.635 ;
        RECT  3.255 1.040 3.335 1.480 ;
        RECT  3.155 0.750 3.220 0.920 ;
        RECT  3.065 0.750 3.155 1.485 ;
        RECT  2.425 1.395 3.065 1.485 ;
        RECT  2.880 0.525 2.975 0.940 ;
        RECT  2.790 1.175 2.900 1.285 ;
        RECT  2.700 0.275 2.790 1.285 ;
        RECT  2.515 0.275 2.610 1.285 ;
        RECT  1.390 0.275 2.515 0.385 ;
        RECT  2.330 0.495 2.425 1.485 ;
        RECT  2.325 0.495 2.330 1.295 ;
        RECT  2.290 1.085 2.325 1.295 ;
        RECT  1.145 1.425 2.240 1.525 ;
        RECT  2.200 0.525 2.225 0.635 ;
        RECT  2.110 0.525 2.200 1.295 ;
        RECT  1.770 0.525 2.110 0.635 ;
        RECT  1.965 1.185 2.110 1.295 ;
        RECT  1.910 0.745 2.020 1.075 ;
        RECT  1.500 0.975 1.910 1.075 ;
        RECT  1.660 0.525 1.770 0.865 ;
        RECT  1.410 0.490 1.500 1.280 ;
        RECT  1.270 0.490 1.410 0.590 ;
        RECT  1.235 1.170 1.410 1.280 ;
        RECT  1.055 1.105 1.145 1.525 ;
        RECT  0.730 1.105 1.055 1.195 ;
        RECT  0.730 0.780 0.830 0.890 ;
        RECT  0.685 0.565 0.730 1.195 ;
        RECT  0.640 0.275 0.685 1.480 ;
        RECT  0.575 0.275 0.640 0.665 ;
        RECT  0.575 1.030 0.640 1.480 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.310 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.185 1.210 0.320 1.310 ;
        RECT  0.075 0.275 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.485 ;
    END
END DFND1

MACRO DFND2
    CLASS CORE ;
    FOREIGN DFND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.575 4.550 1.140 ;
        RECT  4.430 0.575 4.450 0.675 ;
        RECT  4.430 1.040 4.450 1.140 ;
        RECT  4.320 0.275 4.430 0.675 ;
        RECT  4.320 1.040 4.430 1.480 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.515 3.950 1.490 ;
        RECT  3.750 0.515 3.850 0.625 ;
        RECT  3.800 1.040 3.850 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.700 1.300 0.900 ;
        RECT  1.050 0.500 1.150 0.900 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.690 -0.165 4.800 0.165 ;
        RECT  4.580 -0.165 4.690 0.475 ;
        RECT  0.945 -0.165 4.580 0.165 ;
        RECT  0.835 -0.165 0.945 0.670 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.690 1.635 4.800 1.965 ;
        RECT  4.580 1.270 4.690 1.965 ;
        RECT  4.170 1.635 4.580 1.965 ;
        RECT  4.060 1.040 4.170 1.965 ;
        RECT  3.635 1.635 4.060 1.965 ;
        RECT  3.525 1.040 3.635 1.965 ;
        RECT  0.945 1.635 3.525 1.965 ;
        RECT  0.835 1.305 0.945 1.965 ;
        RECT  0.000 1.635 0.835 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.210 0.780 4.340 0.890 ;
        RECT  4.120 0.275 4.210 0.890 ;
        RECT  2.790 0.275 4.120 0.375 ;
        RECT  3.425 0.780 3.760 0.890 ;
        RECT  3.365 0.515 3.425 1.150 ;
        RECT  3.335 0.515 3.365 1.480 ;
        RECT  2.975 0.515 3.335 0.625 ;
        RECT  3.255 1.040 3.335 1.480 ;
        RECT  3.155 0.750 3.220 0.920 ;
        RECT  3.065 0.750 3.155 1.485 ;
        RECT  2.425 1.395 3.065 1.485 ;
        RECT  2.880 0.515 2.975 0.940 ;
        RECT  2.790 1.125 2.900 1.235 ;
        RECT  2.700 0.275 2.790 1.235 ;
        RECT  2.515 0.275 2.610 1.285 ;
        RECT  1.390 0.275 2.515 0.385 ;
        RECT  2.330 0.495 2.425 1.485 ;
        RECT  2.325 0.495 2.330 1.295 ;
        RECT  2.290 1.085 2.325 1.295 ;
        RECT  1.145 1.425 2.240 1.525 ;
        RECT  2.200 0.525 2.225 0.635 ;
        RECT  2.110 0.525 2.200 1.295 ;
        RECT  1.770 0.525 2.110 0.635 ;
        RECT  1.965 1.185 2.110 1.295 ;
        RECT  1.910 0.745 2.020 1.075 ;
        RECT  1.500 0.975 1.910 1.075 ;
        RECT  1.660 0.525 1.770 0.865 ;
        RECT  1.410 0.490 1.500 1.280 ;
        RECT  1.270 0.490 1.410 0.590 ;
        RECT  1.235 1.170 1.410 1.280 ;
        RECT  1.055 1.105 1.145 1.525 ;
        RECT  0.730 1.105 1.055 1.195 ;
        RECT  0.730 0.780 0.830 0.890 ;
        RECT  0.685 0.565 0.730 1.195 ;
        RECT  0.640 0.275 0.685 1.480 ;
        RECT  0.575 0.275 0.640 0.665 ;
        RECT  0.575 1.030 0.640 1.480 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.310 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.185 1.210 0.320 1.310 ;
        RECT  0.075 0.275 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.485 ;
    END
END DFND2

MACRO DFND4
    CLASS CORE ;
    FOREIGN DFND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.275 5.950 0.675 ;
        RECT  5.850 1.040 5.950 1.490 ;
        RECT  5.765 0.275 5.850 1.490 ;
        RECT  5.550 0.505 5.765 1.210 ;
        RECT  5.375 0.505 5.550 0.675 ;
        RECT  5.375 1.040 5.550 1.210 ;
        RECT  5.265 0.275 5.375 0.675 ;
        RECT  5.265 1.040 5.375 1.480 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.515 4.905 0.625 ;
        RECT  4.745 1.040 4.855 1.480 ;
        RECT  4.650 1.040 4.745 1.150 ;
        RECT  4.350 0.515 4.650 1.150 ;
        RECT  4.185 0.515 4.350 0.625 ;
        RECT  4.345 1.040 4.350 1.150 ;
        RECT  4.235 1.040 4.345 1.480 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.700 1.300 0.900 ;
        RECT  1.050 0.500 1.150 0.900 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 6.200 0.165 ;
        RECT  0.835 -0.165 0.945 0.670 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.115 1.635 6.200 1.965 ;
        RECT  5.005 1.040 5.115 1.965 ;
        RECT  4.085 1.635 5.005 1.965 ;
        RECT  3.975 1.040 4.085 1.965 ;
        RECT  0.945 1.635 3.975 1.965 ;
        RECT  0.835 1.305 0.945 1.965 ;
        RECT  0.000 1.635 0.835 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.375 0.505 5.450 0.675 ;
        RECT  5.375 1.040 5.450 1.210 ;
        RECT  5.265 0.275 5.375 0.675 ;
        RECT  5.265 1.040 5.375 1.480 ;
        RECT  4.750 0.515 4.905 0.625 ;
        RECT  4.750 1.040 4.855 1.480 ;
        RECT  4.185 0.515 4.250 0.625 ;
        RECT  4.235 1.040 4.250 1.480 ;
        RECT  5.155 0.780 5.350 0.890 ;
        RECT  5.065 0.315 5.155 0.890 ;
        RECT  2.790 0.315 5.065 0.425 ;
        RECT  3.885 0.780 4.240 0.890 ;
        RECT  3.825 0.515 3.885 1.150 ;
        RECT  3.790 0.515 3.825 1.480 ;
        RECT  3.075 0.515 3.790 0.625 ;
        RECT  3.715 1.040 3.790 1.480 ;
        RECT  3.580 0.780 3.680 0.890 ;
        RECT  3.490 0.780 3.580 1.485 ;
        RECT  2.425 1.395 3.490 1.485 ;
        RECT  2.790 1.125 3.400 1.235 ;
        RECT  2.965 0.515 3.075 0.940 ;
        RECT  2.700 0.315 2.790 1.235 ;
        RECT  2.515 0.275 2.610 1.285 ;
        RECT  1.390 0.275 2.515 0.385 ;
        RECT  2.330 0.495 2.425 1.485 ;
        RECT  2.325 0.495 2.330 1.295 ;
        RECT  2.290 1.085 2.325 1.295 ;
        RECT  1.145 1.425 2.240 1.525 ;
        RECT  2.200 0.525 2.225 0.635 ;
        RECT  2.110 0.525 2.200 1.295 ;
        RECT  1.770 0.525 2.110 0.635 ;
        RECT  1.965 1.185 2.110 1.295 ;
        RECT  1.910 0.745 2.020 1.075 ;
        RECT  1.500 0.975 1.910 1.075 ;
        RECT  1.660 0.525 1.770 0.865 ;
        RECT  1.410 0.490 1.500 1.280 ;
        RECT  1.270 0.490 1.410 0.590 ;
        RECT  1.235 1.170 1.410 1.280 ;
        RECT  1.055 1.105 1.145 1.525 ;
        RECT  0.730 1.105 1.055 1.195 ;
        RECT  0.730 0.780 0.830 0.890 ;
        RECT  0.685 0.565 0.730 1.195 ;
        RECT  0.640 0.275 0.685 1.480 ;
        RECT  0.575 0.275 0.640 0.665 ;
        RECT  0.575 1.030 0.640 1.480 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.310 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.185 1.210 0.320 1.310 ;
        RECT  0.075 0.275 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.485 ;
    END
END DFND4

MACRO DFNSND1
    CLASS CORE ;
    FOREIGN DFNSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0826 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.235 0.710 3.550 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.015 0.525 4.120 1.125 ;
        RECT  3.955 0.525 4.015 0.635 ;
        RECT  3.865 1.015 4.015 1.125 ;
        RECT  3.845 0.310 3.955 0.635 ;
        RECT  3.650 0.310 3.845 0.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.275 4.750 1.490 ;
        RECT  4.615 0.275 4.640 0.650 ;
        RECT  4.615 1.040 4.640 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0486 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.355 0.890 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.265 1.635 4.800 1.965 ;
        RECT  3.095 1.400 3.265 1.965 ;
        RECT  2.400 1.635 3.095 1.965 ;
        RECT  2.210 1.425 2.400 1.965 ;
        RECT  0.000 1.635 2.210 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.505 0.750 4.550 0.920 ;
        RECT  4.415 0.300 4.505 1.505 ;
        RECT  4.065 0.300 4.415 0.415 ;
        RECT  4.080 1.395 4.415 1.505 ;
        RECT  4.210 0.750 4.325 1.305 ;
        RECT  3.990 1.215 4.210 1.305 ;
        RECT  3.455 1.410 4.080 1.505 ;
        RECT  3.890 1.215 3.990 1.310 ;
        RECT  2.810 1.220 3.890 1.310 ;
        RECT  3.770 0.750 3.845 0.920 ;
        RECT  3.680 0.750 3.770 1.130 ;
        RECT  3.115 1.015 3.680 1.130 ;
        RECT  3.115 0.510 3.310 0.620 ;
        RECT  3.015 0.510 3.115 1.130 ;
        RECT  2.650 0.510 3.015 0.655 ;
        RECT  2.920 1.015 3.015 1.130 ;
        RECT  2.670 0.275 2.915 0.390 ;
        RECT  2.700 0.855 2.810 1.310 ;
        RECT  2.535 0.855 2.700 0.945 ;
        RECT  0.430 0.275 2.670 0.370 ;
        RECT  2.495 1.245 2.605 1.525 ;
        RECT  2.265 1.055 2.590 1.155 ;
        RECT  2.420 0.495 2.535 0.945 ;
        RECT  1.695 1.245 2.495 1.335 ;
        RECT  2.175 0.480 2.265 1.155 ;
        RECT  1.695 1.055 2.175 1.155 ;
        RECT  1.825 0.480 1.935 0.920 ;
        RECT  0.960 0.480 1.825 0.590 ;
        RECT  1.605 0.730 1.695 1.155 ;
        RECT  1.605 1.245 1.695 1.465 ;
        RECT  0.780 1.355 1.605 1.465 ;
        RECT  0.960 1.095 1.420 1.205 ;
        RECT  0.870 0.480 0.960 1.205 ;
        RECT  0.670 0.460 0.780 1.465 ;
        RECT  0.540 0.460 0.670 0.580 ;
        RECT  0.575 1.295 0.670 1.465 ;
        RECT  0.430 0.750 0.510 0.920 ;
        RECT  0.320 0.275 0.430 1.310 ;
        RECT  0.185 0.275 0.320 0.370 ;
        RECT  0.185 1.210 0.320 1.310 ;
        RECT  0.075 0.275 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.485 ;
    END
END DFNSND1

MACRO DFNSND2
    CLASS CORE ;
    FOREIGN DFNSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0826 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.750 3.410 0.920 ;
        RECT  3.250 0.510 3.350 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.540 4.150 1.125 ;
        RECT  3.915 0.540 4.050 0.650 ;
        RECT  3.920 1.015 4.050 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.275 5.150 1.490 ;
        RECT  4.965 0.275 5.050 0.655 ;
        RECT  4.965 1.040 5.050 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0416 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.730 1.290 0.900 ;
        RECT  1.050 0.500 1.160 0.900 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 5.400 0.165 ;
        RECT  0.835 -0.165 0.945 0.670 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.325 1.635 5.400 1.965 ;
        RECT  3.145 1.395 3.325 1.965 ;
        RECT  2.435 1.635 3.145 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.945 1.635 2.245 1.965 ;
        RECT  0.835 1.305 0.945 1.965 ;
        RECT  0.000 1.635 0.835 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.855 0.750 4.940 0.920 ;
        RECT  4.765 0.340 4.855 1.505 ;
        RECT  3.640 0.340 4.765 0.450 ;
        RECT  4.435 1.395 4.765 1.505 ;
        RECT  4.465 0.730 4.575 1.305 ;
        RECT  2.845 1.215 4.465 1.305 ;
        RECT  3.820 0.750 3.950 0.920 ;
        RECT  3.730 0.750 3.820 1.125 ;
        RECT  3.150 1.015 3.730 1.125 ;
        RECT  3.530 0.340 3.640 0.920 ;
        RECT  3.150 0.290 3.345 0.400 ;
        RECT  3.055 0.290 3.150 1.125 ;
        RECT  3.050 0.510 3.055 1.125 ;
        RECT  2.685 0.510 3.050 0.655 ;
        RECT  2.955 1.015 3.050 1.125 ;
        RECT  2.705 0.275 2.950 0.390 ;
        RECT  2.735 0.855 2.845 1.305 ;
        RECT  2.570 0.855 2.735 0.945 ;
        RECT  1.350 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.300 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.570 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.210 0.480 2.300 1.155 ;
        RECT  1.730 1.055 2.210 1.155 ;
        RECT  1.860 0.480 1.970 0.920 ;
        RECT  1.540 0.480 1.860 0.590 ;
        RECT  1.640 0.730 1.730 1.155 ;
        RECT  1.640 1.245 1.730 1.465 ;
        RECT  1.155 1.355 1.640 1.465 ;
        RECT  1.430 0.480 1.540 1.205 ;
        RECT  1.250 0.480 1.430 0.590 ;
        RECT  1.245 1.095 1.430 1.205 ;
        RECT  1.055 1.105 1.155 1.465 ;
        RECT  0.730 1.105 1.055 1.195 ;
        RECT  0.730 0.780 0.830 0.890 ;
        RECT  0.685 0.565 0.730 1.195 ;
        RECT  0.640 0.275 0.685 1.480 ;
        RECT  0.575 0.275 0.640 0.665 ;
        RECT  0.575 1.030 0.640 1.480 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.310 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.185 1.210 0.320 1.310 ;
        RECT  0.075 0.275 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.485 ;
    END
END DFNSND2

MACRO DFNSND4
    CLASS CORE ;
    FOREIGN DFNSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1093 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.710 3.450 0.900 ;
        RECT  3.250 0.510 3.350 0.900 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.495 4.625 0.680 ;
        RECT  4.450 1.020 4.610 1.245 ;
        RECT  4.170 0.495 4.450 1.245 ;
        RECT  3.915 0.495 4.170 0.680 ;
        RECT  3.960 1.020 4.170 1.245 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.310 6.150 0.670 ;
        RECT  6.050 1.075 6.150 1.410 ;
        RECT  5.750 0.310 6.050 1.410 ;
        RECT  5.430 0.310 5.750 0.670 ;
        RECT  5.430 1.075 5.750 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0416 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.730 1.290 0.900 ;
        RECT  1.050 0.500 1.160 0.900 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 6.400 0.165 ;
        RECT  0.835 -0.165 0.945 0.670 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.345 1.635 6.400 1.965 ;
        RECT  3.175 1.395 3.345 1.965 ;
        RECT  2.435 1.635 3.175 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.945 1.635 2.245 1.965 ;
        RECT  0.835 1.305 0.945 1.965 ;
        RECT  0.000 1.635 0.835 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.430 0.310 5.650 0.670 ;
        RECT  5.430 1.075 5.650 1.410 ;
        RECT  4.550 0.495 4.625 0.680 ;
        RECT  4.550 1.020 4.610 1.245 ;
        RECT  3.915 0.495 4.050 0.680 ;
        RECT  3.960 1.020 4.050 1.245 ;
        RECT  5.315 0.780 5.615 0.890 ;
        RECT  5.210 0.295 5.315 1.160 ;
        RECT  5.085 0.295 5.210 0.405 ;
        RECT  5.085 1.050 5.210 1.160 ;
        RECT  4.810 0.780 5.100 0.895 ;
        RECT  4.955 0.295 5.085 0.650 ;
        RECT  4.960 1.050 5.085 1.470 ;
        RECT  3.670 0.295 4.955 0.405 ;
        RECT  4.710 0.780 4.810 1.455 ;
        RECT  3.815 1.355 4.710 1.455 ;
        RECT  3.850 0.780 4.060 0.890 ;
        RECT  3.760 0.780 3.850 1.125 ;
        RECT  3.715 1.215 3.815 1.455 ;
        RECT  3.140 1.015 3.760 1.125 ;
        RECT  2.825 1.215 3.715 1.305 ;
        RECT  3.560 0.295 3.670 0.920 ;
        RECT  3.140 0.290 3.335 0.390 ;
        RECT  3.040 0.290 3.140 1.125 ;
        RECT  2.685 0.490 3.040 0.655 ;
        RECT  2.955 1.015 3.040 1.125 ;
        RECT  2.705 0.275 2.950 0.390 ;
        RECT  2.735 0.855 2.825 1.305 ;
        RECT  2.570 0.855 2.735 0.945 ;
        RECT  1.350 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.300 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.570 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.210 0.480 2.300 1.155 ;
        RECT  1.730 1.055 2.210 1.155 ;
        RECT  1.860 0.480 1.970 0.920 ;
        RECT  1.540 0.480 1.860 0.590 ;
        RECT  1.640 0.730 1.730 1.155 ;
        RECT  1.640 1.245 1.730 1.465 ;
        RECT  1.155 1.355 1.640 1.465 ;
        RECT  1.430 0.480 1.540 1.205 ;
        RECT  1.250 0.480 1.430 0.590 ;
        RECT  1.245 1.095 1.430 1.205 ;
        RECT  1.055 1.105 1.155 1.465 ;
        RECT  0.730 1.105 1.055 1.195 ;
        RECT  0.730 0.780 0.830 0.890 ;
        RECT  0.685 0.565 0.730 1.195 ;
        RECT  0.640 0.275 0.685 1.480 ;
        RECT  0.575 0.275 0.640 0.665 ;
        RECT  0.575 1.030 0.640 1.480 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.310 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.185 1.210 0.320 1.310 ;
        RECT  0.075 0.275 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.485 ;
    END
END DFNSND4

MACRO DFQD1
    CLASS CORE ;
    FOREIGN DFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.595 0.290 3.750 1.500 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.710 1.260 0.920 ;
        RECT  1.050 0.710 1.170 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.670 0.155 1.110 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.915 -0.165 3.800 0.165 ;
        RECT  2.745 -0.165 2.915 0.470 ;
        RECT  0.935 -0.165 2.745 0.165 ;
        RECT  0.760 -0.165 0.935 0.395 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.930 1.635 3.800 1.965 ;
        RECT  2.775 1.450 2.930 1.965 ;
        RECT  0.000 1.635 2.775 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.350 0.570 3.480 1.420 ;
        RECT  3.190 0.570 3.350 0.660 ;
        RECT  3.040 1.315 3.350 1.420 ;
        RECT  3.080 0.285 3.190 0.660 ;
        RECT  2.985 0.750 3.095 1.220 ;
        RECT  2.860 0.570 3.080 0.660 ;
        RECT  2.320 1.120 2.985 1.220 ;
        RECT  2.750 0.570 2.860 0.920 ;
        RECT  2.500 0.865 2.645 0.995 ;
        RECT  2.410 0.275 2.500 0.995 ;
        RECT  0.420 1.430 2.440 1.525 ;
        RECT  2.285 0.275 2.410 0.365 ;
        RECT  2.210 0.455 2.320 1.220 ;
        RECT  2.115 0.255 2.285 0.365 ;
        RECT  2.010 0.475 2.120 1.340 ;
        RECT  1.125 0.275 2.115 0.365 ;
        RECT  1.715 0.475 2.010 0.600 ;
        RECT  1.830 0.750 1.920 1.315 ;
        RECT  1.500 1.205 1.830 1.315 ;
        RECT  1.600 0.475 1.715 0.920 ;
        RECT  1.390 0.480 1.500 1.315 ;
        RECT  1.215 0.480 1.390 0.605 ;
        RECT  1.205 1.205 1.390 1.315 ;
        RECT  1.025 0.275 1.125 0.620 ;
        RECT  0.800 0.500 1.025 0.620 ;
        RECT  0.680 0.500 0.800 1.160 ;
        RECT  0.540 0.500 0.680 0.660 ;
        RECT  0.525 1.040 0.680 1.160 ;
        RECT  0.420 0.770 0.570 0.900 ;
        RECT  0.320 0.460 0.420 1.525 ;
        RECT  0.180 0.460 0.320 0.560 ;
        RECT  0.075 1.230 0.320 1.400 ;
        RECT  0.080 0.370 0.180 0.560 ;
    END
END DFQD1

MACRO DFQD2
    CLASS CORE ;
    FOREIGN DFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.565 0.290 3.750 1.500 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.710 1.260 0.920 ;
        RECT  1.050 0.710 1.170 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.670 0.155 1.110 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.915 -0.165 4.000 0.165 ;
        RECT  2.745 -0.165 2.915 0.470 ;
        RECT  0.935 -0.165 2.745 0.165 ;
        RECT  0.760 -0.165 0.935 0.395 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.930 1.635 4.000 1.965 ;
        RECT  2.775 1.450 2.930 1.965 ;
        RECT  0.000 1.635 2.775 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.345 0.570 3.455 1.420 ;
        RECT  3.190 0.570 3.345 0.660 ;
        RECT  3.040 1.315 3.345 1.420 ;
        RECT  3.080 0.285 3.190 0.660 ;
        RECT  2.985 0.750 3.095 1.220 ;
        RECT  2.860 0.570 3.080 0.660 ;
        RECT  2.320 1.120 2.985 1.220 ;
        RECT  2.750 0.570 2.860 0.920 ;
        RECT  2.500 0.865 2.645 0.995 ;
        RECT  2.410 0.275 2.500 0.995 ;
        RECT  0.420 1.430 2.440 1.525 ;
        RECT  2.285 0.275 2.410 0.365 ;
        RECT  2.210 0.455 2.320 1.220 ;
        RECT  2.115 0.255 2.285 0.365 ;
        RECT  2.010 0.475 2.120 1.340 ;
        RECT  1.125 0.275 2.115 0.365 ;
        RECT  1.715 0.475 2.010 0.600 ;
        RECT  1.830 0.750 1.920 1.315 ;
        RECT  1.500 1.205 1.830 1.315 ;
        RECT  1.600 0.475 1.715 0.920 ;
        RECT  1.390 0.480 1.500 1.315 ;
        RECT  1.215 0.480 1.390 0.605 ;
        RECT  1.205 1.205 1.390 1.315 ;
        RECT  1.025 0.275 1.125 0.620 ;
        RECT  0.800 0.500 1.025 0.620 ;
        RECT  0.680 0.500 0.800 1.160 ;
        RECT  0.540 0.500 0.680 0.660 ;
        RECT  0.525 1.040 0.680 1.160 ;
        RECT  0.420 0.770 0.570 0.900 ;
        RECT  0.320 0.460 0.420 1.525 ;
        RECT  0.180 0.460 0.320 0.560 ;
        RECT  0.075 1.230 0.320 1.400 ;
        RECT  0.080 0.370 0.180 0.560 ;
    END
END DFQD2

MACRO DFQD4
    CLASS CORE ;
    FOREIGN DFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.110 0.290 4.240 0.695 ;
        RECT  4.110 1.005 4.240 1.500 ;
        RECT  4.050 0.530 4.110 0.695 ;
        RECT  4.050 1.005 4.110 1.215 ;
        RECT  3.750 0.530 4.050 1.215 ;
        RECT  3.720 0.530 3.750 0.695 ;
        RECT  3.720 1.005 3.750 1.215 ;
        RECT  3.590 0.290 3.720 0.695 ;
        RECT  3.585 1.005 3.720 1.500 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.710 1.260 0.920 ;
        RECT  1.050 0.710 1.170 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.770 0.200 0.960 ;
        RECT  0.045 0.670 0.155 1.110 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.490 -0.165 4.600 0.165 ;
        RECT  4.380 -0.165 4.490 0.705 ;
        RECT  4.000 -0.165 4.380 0.165 ;
        RECT  3.830 -0.165 4.000 0.420 ;
        RECT  3.450 -0.165 3.830 0.165 ;
        RECT  3.340 -0.165 3.450 0.465 ;
        RECT  2.915 -0.165 3.340 0.165 ;
        RECT  2.745 -0.165 2.915 0.470 ;
        RECT  0.935 -0.165 2.745 0.165 ;
        RECT  0.760 -0.165 0.935 0.395 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.490 1.635 4.600 1.965 ;
        RECT  4.380 1.040 4.490 1.965 ;
        RECT  3.970 1.635 4.380 1.965 ;
        RECT  3.860 1.325 3.970 1.965 ;
        RECT  2.930 1.635 3.860 1.965 ;
        RECT  2.775 1.450 2.930 1.965 ;
        RECT  0.000 1.635 2.775 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.150 0.290 4.240 0.695 ;
        RECT  4.150 1.005 4.240 1.500 ;
        RECT  3.590 0.290 3.650 0.695 ;
        RECT  3.585 1.005 3.650 1.500 ;
        RECT  3.405 0.785 3.595 0.895 ;
        RECT  3.295 0.570 3.405 1.450 ;
        RECT  3.190 0.570 3.295 0.660 ;
        RECT  3.040 1.335 3.295 1.450 ;
        RECT  3.080 0.285 3.190 0.660 ;
        RECT  2.985 0.750 3.095 1.220 ;
        RECT  2.860 0.570 3.080 0.660 ;
        RECT  2.320 1.120 2.985 1.220 ;
        RECT  2.750 0.570 2.860 0.920 ;
        RECT  2.500 0.865 2.645 0.995 ;
        RECT  2.410 0.275 2.500 0.995 ;
        RECT  0.420 1.430 2.440 1.525 ;
        RECT  2.285 0.275 2.410 0.365 ;
        RECT  2.210 0.455 2.320 1.220 ;
        RECT  2.115 0.255 2.285 0.365 ;
        RECT  2.010 0.475 2.120 1.340 ;
        RECT  1.125 0.275 2.115 0.365 ;
        RECT  1.715 0.475 2.010 0.600 ;
        RECT  1.830 0.750 1.920 1.315 ;
        RECT  1.500 1.205 1.830 1.315 ;
        RECT  1.600 0.475 1.715 0.920 ;
        RECT  1.390 0.480 1.500 1.315 ;
        RECT  1.215 0.480 1.390 0.605 ;
        RECT  1.205 1.205 1.390 1.315 ;
        RECT  1.025 0.275 1.125 0.620 ;
        RECT  0.800 0.500 1.025 0.620 ;
        RECT  0.680 0.500 0.800 1.160 ;
        RECT  0.540 0.500 0.680 0.660 ;
        RECT  0.525 1.040 0.680 1.160 ;
        RECT  0.420 0.770 0.570 0.900 ;
        RECT  0.320 0.460 0.420 1.525 ;
        RECT  0.180 0.460 0.320 0.560 ;
        RECT  0.075 1.230 0.320 1.400 ;
        RECT  0.080 0.370 0.180 0.560 ;
    END
END DFQD4

MACRO DFSND1
    CLASS CORE ;
    FOREIGN DFSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0823 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 0.750 3.410 0.920 ;
        RECT  3.250 0.510 3.370 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.510 4.155 1.125 ;
        RECT  3.935 0.510 4.050 0.620 ;
        RECT  3.965 1.015 4.050 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.275 4.950 1.480 ;
        RECT  4.755 0.275 4.850 0.680 ;
        RECT  4.755 1.040 4.850 1.480 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.290 0.930 ;
        RECT  1.050 0.760 1.150 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 5.000 0.165 ;
        RECT  0.835 -0.165 0.945 0.450 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.890 1.635 5.000 1.965 ;
        RECT  3.720 1.395 3.890 1.965 ;
        RECT  3.325 1.635 3.720 1.965 ;
        RECT  3.145 1.395 3.325 1.965 ;
        RECT  2.435 1.635 3.145 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.000 1.635 2.245 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.645 0.780 4.760 0.890 ;
        RECT  4.555 0.310 4.645 1.505 ;
        RECT  3.640 0.310 4.555 0.420 ;
        RECT  4.185 1.395 4.555 1.505 ;
        RECT  4.310 0.730 4.425 1.305 ;
        RECT  2.845 1.215 4.310 1.305 ;
        RECT  3.845 0.780 3.960 0.890 ;
        RECT  3.745 0.780 3.845 1.125 ;
        RECT  3.160 1.015 3.745 1.125 ;
        RECT  3.530 0.310 3.640 0.920 ;
        RECT  3.160 0.305 3.345 0.415 ;
        RECT  3.070 0.305 3.160 1.125 ;
        RECT  2.700 0.510 3.070 0.655 ;
        RECT  2.955 1.015 3.070 1.125 ;
        RECT  2.705 0.275 2.980 0.390 ;
        RECT  2.735 0.855 2.845 1.305 ;
        RECT  2.580 0.855 2.735 0.945 ;
        RECT  1.170 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.335 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.580 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.220 0.480 2.335 1.155 ;
        RECT  1.755 1.055 2.220 1.155 ;
        RECT  1.885 0.480 1.995 0.920 ;
        RECT  1.540 0.480 1.885 0.590 ;
        RECT  1.665 0.730 1.755 1.155 ;
        RECT  1.640 1.245 1.730 1.470 ;
        RECT  0.430 1.380 1.640 1.470 ;
        RECT  1.430 0.480 1.540 1.250 ;
        RECT  1.270 0.480 1.430 0.590 ;
        RECT  1.260 1.140 1.430 1.250 ;
        RECT  1.080 0.275 1.170 0.655 ;
        RECT  0.840 0.560 1.080 0.655 ;
        RECT  0.750 0.560 0.840 1.265 ;
        RECT  0.685 0.560 0.750 0.655 ;
        RECT  0.535 1.130 0.750 1.265 ;
        RECT  0.575 0.275 0.685 0.655 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.470 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.075 1.300 0.320 1.470 ;
        RECT  0.075 0.275 0.185 0.590 ;
    END
END DFSND1

MACRO DFSND2
    CLASS CORE ;
    FOREIGN DFSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0823 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 0.750 3.410 0.920 ;
        RECT  3.250 0.510 3.370 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.540 4.150 1.125 ;
        RECT  3.915 0.540 4.050 0.650 ;
        RECT  3.920 1.015 4.050 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.275 5.150 1.490 ;
        RECT  4.965 0.275 5.050 0.650 ;
        RECT  4.965 1.040 5.050 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.290 0.930 ;
        RECT  1.050 0.760 1.150 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 5.400 0.165 ;
        RECT  0.835 -0.165 0.945 0.450 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.325 1.635 5.400 1.965 ;
        RECT  3.145 1.395 3.325 1.965 ;
        RECT  2.435 1.635 3.145 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.000 1.635 2.245 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.855 0.750 4.940 0.920 ;
        RECT  4.765 0.340 4.855 1.505 ;
        RECT  3.640 0.340 4.765 0.450 ;
        RECT  4.435 1.395 4.765 1.505 ;
        RECT  4.465 0.730 4.575 1.305 ;
        RECT  2.845 1.215 4.465 1.305 ;
        RECT  3.820 0.750 3.940 0.920 ;
        RECT  3.730 0.750 3.820 1.125 ;
        RECT  3.160 1.015 3.730 1.125 ;
        RECT  3.530 0.340 3.640 0.920 ;
        RECT  3.160 0.305 3.345 0.415 ;
        RECT  3.070 0.305 3.160 1.125 ;
        RECT  2.700 0.510 3.070 0.655 ;
        RECT  2.955 1.015 3.070 1.125 ;
        RECT  2.705 0.275 2.980 0.390 ;
        RECT  2.735 0.855 2.845 1.305 ;
        RECT  2.580 0.855 2.735 0.945 ;
        RECT  1.170 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.335 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.580 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.220 0.480 2.335 1.155 ;
        RECT  1.755 1.055 2.220 1.155 ;
        RECT  1.885 0.480 1.995 0.920 ;
        RECT  1.540 0.480 1.885 0.590 ;
        RECT  1.665 0.730 1.755 1.155 ;
        RECT  1.640 1.245 1.730 1.470 ;
        RECT  0.430 1.380 1.640 1.470 ;
        RECT  1.430 0.480 1.540 1.250 ;
        RECT  1.270 0.480 1.430 0.590 ;
        RECT  1.260 1.140 1.430 1.250 ;
        RECT  1.080 0.275 1.170 0.655 ;
        RECT  0.840 0.560 1.080 0.655 ;
        RECT  0.750 0.560 0.840 1.265 ;
        RECT  0.685 0.560 0.750 0.655 ;
        RECT  0.535 1.130 0.750 1.265 ;
        RECT  0.575 0.275 0.685 0.655 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.470 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.075 1.300 0.320 1.470 ;
        RECT  0.075 0.275 0.185 0.590 ;
    END
END DFSND2

MACRO DFSND4
    CLASS CORE ;
    FOREIGN DFSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1093 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.710 3.450 0.900 ;
        RECT  3.250 0.510 3.350 0.900 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.495 4.625 0.680 ;
        RECT  4.450 1.020 4.610 1.245 ;
        RECT  4.170 0.495 4.450 1.245 ;
        RECT  3.915 0.495 4.170 0.680 ;
        RECT  3.960 1.020 4.170 1.245 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.310 6.150 0.680 ;
        RECT  6.050 1.060 6.150 1.430 ;
        RECT  5.750 0.310 6.050 1.430 ;
        RECT  5.465 0.310 5.750 0.680 ;
        RECT  5.465 1.060 5.750 1.430 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.290 0.930 ;
        RECT  1.050 0.760 1.150 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 6.400 0.165 ;
        RECT  0.835 -0.165 0.945 0.450 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.345 1.635 6.400 1.965 ;
        RECT  3.175 1.395 3.345 1.965 ;
        RECT  2.435 1.635 3.175 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.000 1.635 2.245 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.465 0.310 5.650 0.680 ;
        RECT  5.465 1.060 5.650 1.430 ;
        RECT  4.550 0.495 4.625 0.680 ;
        RECT  4.550 1.020 4.610 1.245 ;
        RECT  3.915 0.495 4.050 0.680 ;
        RECT  3.960 1.020 4.050 1.245 ;
        RECT  5.315 0.780 5.615 0.890 ;
        RECT  5.210 0.295 5.315 1.160 ;
        RECT  5.085 0.295 5.210 0.405 ;
        RECT  5.085 1.050 5.210 1.160 ;
        RECT  4.810 0.780 5.100 0.895 ;
        RECT  4.955 0.295 5.085 0.650 ;
        RECT  4.960 1.050 5.085 1.470 ;
        RECT  3.670 0.295 4.955 0.405 ;
        RECT  4.710 0.780 4.810 1.455 ;
        RECT  3.815 1.355 4.710 1.455 ;
        RECT  3.850 0.780 4.060 0.890 ;
        RECT  3.760 0.780 3.850 1.125 ;
        RECT  3.715 1.215 3.815 1.455 ;
        RECT  3.160 1.015 3.760 1.125 ;
        RECT  2.845 1.215 3.715 1.305 ;
        RECT  3.560 0.295 3.670 0.920 ;
        RECT  3.160 0.290 3.335 0.390 ;
        RECT  3.070 0.290 3.160 1.125 ;
        RECT  2.700 0.510 3.070 0.655 ;
        RECT  2.955 1.015 3.070 1.125 ;
        RECT  2.705 0.275 2.980 0.390 ;
        RECT  2.735 0.855 2.845 1.305 ;
        RECT  2.580 0.855 2.735 0.945 ;
        RECT  1.170 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.335 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.580 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.220 0.480 2.335 1.155 ;
        RECT  1.755 1.055 2.220 1.155 ;
        RECT  1.885 0.480 1.995 0.920 ;
        RECT  1.540 0.480 1.885 0.590 ;
        RECT  1.665 0.730 1.755 1.155 ;
        RECT  1.640 1.245 1.730 1.470 ;
        RECT  0.430 1.380 1.640 1.470 ;
        RECT  1.430 0.480 1.540 1.250 ;
        RECT  1.270 0.480 1.430 0.590 ;
        RECT  1.260 1.140 1.430 1.250 ;
        RECT  1.080 0.275 1.170 0.655 ;
        RECT  0.840 0.560 1.080 0.655 ;
        RECT  0.750 0.560 0.840 1.265 ;
        RECT  0.685 0.560 0.750 0.655 ;
        RECT  0.535 1.130 0.750 1.265 ;
        RECT  0.575 0.275 0.685 0.655 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.470 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.075 1.300 0.320 1.470 ;
        RECT  0.075 0.275 0.185 0.590 ;
    END
END DFSND4

MACRO DFSNQD1
    CLASS CORE ;
    FOREIGN DFSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0730 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 0.750 3.410 0.920 ;
        RECT  3.250 0.510 3.360 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.275 4.550 1.490 ;
        RECT  4.415 0.275 4.450 0.650 ;
        RECT  4.415 1.040 4.450 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.290 0.930 ;
        RECT  1.050 0.760 1.150 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 4.600 0.165 ;
        RECT  0.835 -0.165 0.945 0.450 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.300 1.635 4.600 1.965 ;
        RECT  3.120 1.415 3.300 1.965 ;
        RECT  2.435 1.635 3.120 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.000 1.635 2.245 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.750 4.360 0.920 ;
        RECT  4.215 0.310 4.305 1.505 ;
        RECT  3.625 0.310 4.215 0.420 ;
        RECT  3.865 1.395 4.215 1.505 ;
        RECT  3.990 0.730 4.105 1.305 ;
        RECT  3.770 1.215 3.990 1.305 ;
        RECT  3.680 1.215 3.770 1.325 ;
        RECT  2.845 1.235 3.680 1.325 ;
        RECT  3.515 0.310 3.625 0.920 ;
        RECT  3.145 1.015 3.590 1.135 ;
        RECT  3.145 0.305 3.330 0.415 ;
        RECT  3.055 0.305 3.145 1.135 ;
        RECT  2.700 0.510 3.055 0.655 ;
        RECT  2.955 1.015 3.055 1.135 ;
        RECT  2.705 0.275 2.955 0.390 ;
        RECT  2.735 0.855 2.845 1.325 ;
        RECT  2.580 0.855 2.735 0.945 ;
        RECT  1.170 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.335 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.580 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.220 0.480 2.335 1.155 ;
        RECT  1.755 1.055 2.220 1.155 ;
        RECT  1.885 0.480 1.995 0.920 ;
        RECT  1.540 0.480 1.885 0.590 ;
        RECT  1.665 0.730 1.755 1.155 ;
        RECT  1.640 1.245 1.730 1.470 ;
        RECT  0.430 1.380 1.640 1.470 ;
        RECT  1.430 0.480 1.540 1.250 ;
        RECT  1.270 0.480 1.430 0.590 ;
        RECT  1.260 1.140 1.430 1.250 ;
        RECT  1.080 0.275 1.170 0.655 ;
        RECT  0.840 0.560 1.080 0.655 ;
        RECT  0.750 0.560 0.840 1.265 ;
        RECT  0.685 0.560 0.750 0.655 ;
        RECT  0.535 1.130 0.750 1.265 ;
        RECT  0.575 0.275 0.685 0.655 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.470 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.075 1.300 0.320 1.470 ;
        RECT  0.075 0.275 0.185 0.590 ;
    END
END DFSNQD1

MACRO DFSNQD2
    CLASS CORE ;
    FOREIGN DFSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0730 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 0.750 3.410 0.920 ;
        RECT  3.250 0.510 3.370 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.580 4.750 1.140 ;
        RECT  4.635 0.580 4.650 0.680 ;
        RECT  4.635 1.040 4.650 1.140 ;
        RECT  4.525 0.275 4.635 0.680 ;
        RECT  4.525 1.040 4.635 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.290 0.930 ;
        RECT  1.050 0.760 1.150 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.910 -0.165 5.000 0.165 ;
        RECT  4.775 -0.165 4.910 0.465 ;
        RECT  4.400 -0.165 4.775 0.165 ;
        RECT  4.230 -0.165 4.400 0.405 ;
        RECT  3.870 -0.165 4.230 0.165 ;
        RECT  3.700 -0.165 3.870 0.405 ;
        RECT  0.945 -0.165 3.700 0.165 ;
        RECT  0.835 -0.165 0.945 0.450 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.915 1.635 5.000 1.965 ;
        RECT  4.775 1.295 4.915 1.965 ;
        RECT  3.875 1.635 4.775 1.965 ;
        RECT  3.705 1.395 3.875 1.965 ;
        RECT  3.325 1.635 3.705 1.965 ;
        RECT  3.145 1.395 3.325 1.965 ;
        RECT  2.435 1.635 3.145 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.000 1.635 2.245 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.365 0.780 4.530 0.890 ;
        RECT  4.255 0.505 4.365 1.505 ;
        RECT  3.640 0.505 4.255 0.615 ;
        RECT  3.965 1.395 4.255 1.505 ;
        RECT  3.995 0.730 4.105 1.305 ;
        RECT  2.845 1.215 3.995 1.305 ;
        RECT  3.530 0.505 3.640 0.920 ;
        RECT  3.160 1.015 3.630 1.125 ;
        RECT  3.160 0.305 3.345 0.415 ;
        RECT  3.070 0.305 3.160 1.125 ;
        RECT  2.700 0.510 3.070 0.655 ;
        RECT  2.955 1.015 3.070 1.125 ;
        RECT  2.705 0.275 2.980 0.390 ;
        RECT  2.735 0.855 2.845 1.305 ;
        RECT  2.580 0.855 2.735 0.945 ;
        RECT  1.170 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.335 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.580 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.220 0.480 2.335 1.155 ;
        RECT  1.755 1.055 2.220 1.155 ;
        RECT  1.885 0.480 1.995 0.920 ;
        RECT  1.540 0.480 1.885 0.590 ;
        RECT  1.665 0.730 1.755 1.155 ;
        RECT  1.640 1.245 1.730 1.470 ;
        RECT  0.430 1.380 1.640 1.470 ;
        RECT  1.430 0.480 1.540 1.250 ;
        RECT  1.270 0.480 1.430 0.590 ;
        RECT  1.260 1.140 1.430 1.250 ;
        RECT  1.080 0.275 1.170 0.655 ;
        RECT  0.840 0.560 1.080 0.655 ;
        RECT  0.750 0.560 0.840 1.265 ;
        RECT  0.685 0.560 0.750 0.655 ;
        RECT  0.535 1.130 0.750 1.265 ;
        RECT  0.575 0.275 0.685 0.655 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.470 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.075 1.300 0.320 1.470 ;
        RECT  0.075 0.275 0.185 0.590 ;
    END
END DFSNQD2

MACRO DFSNQD4
    CLASS CORE ;
    FOREIGN DFSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0730 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 0.710 3.450 0.900 ;
        RECT  3.250 0.510 3.370 0.900 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.310 5.150 0.680 ;
        RECT  5.050 1.060 5.150 1.430 ;
        RECT  4.750 0.310 5.050 1.430 ;
        RECT  4.465 0.310 4.750 0.680 ;
        RECT  4.465 1.060 4.750 1.430 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.760 1.290 0.930 ;
        RECT  1.050 0.760 1.150 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.165 5.400 0.165 ;
        RECT  0.835 -0.165 0.945 0.450 ;
        RECT  0.000 -0.165 0.835 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.635 5.400 1.965 ;
        RECT  3.150 1.395 3.320 1.965 ;
        RECT  2.435 1.635 3.150 1.965 ;
        RECT  2.245 1.425 2.435 1.965 ;
        RECT  0.000 1.635 2.245 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.465 0.310 4.650 0.680 ;
        RECT  4.465 1.060 4.650 1.430 ;
        RECT  4.315 0.780 4.615 0.890 ;
        RECT  4.210 0.295 4.315 1.160 ;
        RECT  4.085 0.295 4.210 0.405 ;
        RECT  4.085 1.050 4.210 1.160 ;
        RECT  3.860 0.780 4.100 0.895 ;
        RECT  3.955 0.295 4.085 0.650 ;
        RECT  3.960 1.050 4.085 1.470 ;
        RECT  3.670 0.295 3.955 0.405 ;
        RECT  3.760 0.780 3.860 1.305 ;
        RECT  2.845 1.215 3.760 1.305 ;
        RECT  3.560 0.295 3.670 0.920 ;
        RECT  3.160 1.015 3.620 1.125 ;
        RECT  3.160 0.305 3.335 0.415 ;
        RECT  3.070 0.305 3.160 1.125 ;
        RECT  2.700 0.510 3.070 0.655 ;
        RECT  2.955 1.015 3.070 1.125 ;
        RECT  2.705 0.275 2.980 0.390 ;
        RECT  2.735 0.855 2.845 1.305 ;
        RECT  2.580 0.855 2.735 0.945 ;
        RECT  1.170 0.275 2.705 0.370 ;
        RECT  2.530 1.245 2.640 1.525 ;
        RECT  2.335 1.055 2.625 1.155 ;
        RECT  2.455 0.495 2.580 0.945 ;
        RECT  1.730 1.245 2.530 1.335 ;
        RECT  2.220 0.480 2.335 1.155 ;
        RECT  1.755 1.055 2.220 1.155 ;
        RECT  1.885 0.480 1.995 0.920 ;
        RECT  1.540 0.480 1.885 0.590 ;
        RECT  1.665 0.730 1.755 1.155 ;
        RECT  1.640 1.245 1.730 1.470 ;
        RECT  0.430 1.380 1.640 1.470 ;
        RECT  1.430 0.480 1.540 1.250 ;
        RECT  1.270 0.480 1.430 0.590 ;
        RECT  1.260 1.140 1.430 1.250 ;
        RECT  1.080 0.275 1.170 0.655 ;
        RECT  0.840 0.560 1.080 0.655 ;
        RECT  0.750 0.560 0.840 1.265 ;
        RECT  0.685 0.560 0.750 0.655 ;
        RECT  0.535 1.130 0.750 1.265 ;
        RECT  0.575 0.275 0.685 0.655 ;
        RECT  0.430 0.750 0.530 0.920 ;
        RECT  0.320 0.490 0.430 1.470 ;
        RECT  0.185 0.490 0.320 0.590 ;
        RECT  0.075 1.300 0.320 1.470 ;
        RECT  0.075 0.275 0.185 0.590 ;
    END
END DFSNQD4

MACRO DFXD1
    CLASS CORE ;
    FOREIGN DFXD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.275 5.350 1.490 ;
        RECT  5.220 0.275 5.250 0.675 ;
        RECT  5.215 1.040 5.250 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.475 4.950 1.140 ;
        RECT  4.725 0.475 4.850 0.675 ;
        RECT  4.835 1.040 4.850 1.140 ;
        RECT  4.725 1.040 4.835 1.490 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        RECT  1.315 0.750 1.445 0.920 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.590 1.100 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.700 1.755 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.480 -0.165 5.400 0.165 ;
        RECT  0.305 -0.165 0.480 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.200 1.635 5.400 1.965 ;
        RECT  3.030 1.195 3.200 1.965 ;
        RECT  0.475 1.635 3.030 1.965 ;
        RECT  0.305 1.415 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.130 0.750 5.160 0.920 ;
        RECT  5.040 0.295 5.130 0.920 ;
        RECT  4.045 0.295 5.040 0.385 ;
        RECT  4.635 0.780 4.760 0.890 ;
        RECT  4.570 0.495 4.635 1.330 ;
        RECT  4.545 0.495 4.570 1.490 ;
        RECT  4.225 0.495 4.545 0.605 ;
        RECT  4.460 1.230 4.545 1.490 ;
        RECT  4.405 0.750 4.455 0.920 ;
        RECT  4.315 0.750 4.405 1.120 ;
        RECT  4.300 1.030 4.315 1.120 ;
        RECT  4.210 1.030 4.300 1.515 ;
        RECT  4.135 0.495 4.225 0.920 ;
        RECT  3.645 1.400 4.210 1.515 ;
        RECT  3.955 0.295 4.045 1.245 ;
        RECT  3.770 0.275 3.860 1.310 ;
        RECT  3.610 0.275 3.770 0.365 ;
        RECT  3.740 0.730 3.770 1.310 ;
        RECT  3.645 0.455 3.680 0.640 ;
        RECT  3.555 0.455 3.645 1.515 ;
        RECT  3.440 0.255 3.610 0.365 ;
        RECT  3.375 0.475 3.465 1.330 ;
        RECT  2.690 0.275 3.440 0.365 ;
        RECT  3.065 0.475 3.375 0.585 ;
        RECT  3.290 1.205 3.375 1.330 ;
        RECT  3.185 0.765 3.285 1.085 ;
        RECT  2.830 0.995 3.185 1.085 ;
        RECT  2.945 0.475 3.065 0.905 ;
        RECT  2.720 0.470 2.830 1.320 ;
        RECT  2.560 0.470 2.720 0.595 ;
        RECT  2.560 1.195 2.720 1.320 ;
        RECT  2.260 0.255 2.470 0.375 ;
        RECT  2.350 0.535 2.460 1.195 ;
        RECT  0.930 1.390 2.450 1.500 ;
        RECT  2.050 0.535 2.350 0.645 ;
        RECT  2.050 1.085 2.350 1.195 ;
        RECT  1.150 0.275 2.260 0.375 ;
        RECT  1.935 0.790 2.170 0.900 ;
        RECT  1.845 0.480 1.935 1.300 ;
        RECT  1.550 0.480 1.845 0.590 ;
        RECT  1.550 1.210 1.845 1.300 ;
        RECT  1.135 0.520 1.300 0.630 ;
        RECT  1.135 1.170 1.220 1.280 ;
        RECT  1.050 0.275 1.150 0.410 ;
        RECT  1.045 0.520 1.135 1.280 ;
        RECT  0.830 0.310 1.050 0.410 ;
        RECT  0.815 1.110 0.930 1.500 ;
        RECT  0.695 0.500 0.805 0.965 ;
        RECT  0.350 0.500 0.695 0.590 ;
        RECT  0.260 0.500 0.350 1.320 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.230 0.260 1.320 ;
        RECT  0.075 0.300 0.185 0.590 ;
        RECT  0.075 1.230 0.185 1.495 ;
    END
END DFXD1

MACRO DFXD2
    CLASS CORE ;
    FOREIGN DFXD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.575 5.950 1.140 ;
        RECT  5.805 0.575 5.850 0.675 ;
        RECT  5.805 1.040 5.850 1.140 ;
        RECT  5.695 0.275 5.805 0.675 ;
        RECT  5.650 1.040 5.805 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.285 0.495 5.350 1.140 ;
        RECT  5.250 0.495 5.285 1.470 ;
        RECT  5.125 0.495 5.250 0.605 ;
        RECT  5.175 1.040 5.250 1.470 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        RECT  1.315 0.750 1.445 0.920 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.590 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.700 1.755 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.065 -0.165 6.200 0.165 ;
        RECT  5.955 -0.165 6.065 0.475 ;
        RECT  3.265 -0.165 5.955 0.165 ;
        RECT  3.095 -0.165 3.265 0.295 ;
        RECT  0.480 -0.165 3.095 0.165 ;
        RECT  0.305 -0.165 0.480 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.065 1.635 6.200 1.965 ;
        RECT  5.955 1.260 6.065 1.965 ;
        RECT  5.545 1.635 5.955 1.965 ;
        RECT  5.435 1.260 5.545 1.965 ;
        RECT  5.025 1.635 5.435 1.965 ;
        RECT  4.915 1.040 5.025 1.965 ;
        RECT  3.200 1.635 4.915 1.965 ;
        RECT  3.200 1.195 3.320 1.305 ;
        RECT  3.085 1.195 3.200 1.965 ;
        RECT  0.500 1.635 3.085 1.965 ;
        RECT  0.330 1.415 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.585 0.780 5.760 0.890 ;
        RECT  5.495 0.295 5.585 0.890 ;
        RECT  4.200 0.295 5.495 0.385 ;
        RECT  4.825 0.775 5.160 0.895 ;
        RECT  4.765 0.495 4.825 1.140 ;
        RECT  4.730 0.495 4.765 1.470 ;
        RECT  4.385 0.495 4.730 0.605 ;
        RECT  4.655 1.040 4.730 1.470 ;
        RECT  4.565 0.750 4.635 0.920 ;
        RECT  4.475 0.750 4.565 1.525 ;
        RECT  3.810 1.435 4.475 1.525 ;
        RECT  4.290 0.495 4.385 0.940 ;
        RECT  4.200 1.035 4.230 1.245 ;
        RECT  4.100 0.295 4.200 1.245 ;
        RECT  4.000 0.275 4.010 1.030 ;
        RECT  3.910 0.275 4.000 1.245 ;
        RECT  3.570 0.275 3.910 0.365 ;
        RECT  3.900 0.930 3.910 1.245 ;
        RECT  3.810 0.455 3.820 0.820 ;
        RECT  3.710 0.455 3.810 1.525 ;
        RECT  3.700 0.710 3.710 1.525 ;
        RECT  3.480 0.275 3.570 0.475 ;
        RECT  3.455 0.565 3.555 1.255 ;
        RECT  2.935 0.385 3.480 0.475 ;
        RECT  3.105 0.565 3.455 0.665 ;
        RECT  3.255 0.765 3.365 1.105 ;
        RECT  2.765 1.015 3.255 1.105 ;
        RECT  2.995 0.565 3.105 0.925 ;
        RECT  2.825 0.275 2.935 0.475 ;
        RECT  2.715 1.015 2.765 1.340 ;
        RECT  2.655 0.415 2.715 1.340 ;
        RECT  2.615 0.415 2.655 1.105 ;
        RECT  0.995 1.390 2.520 1.500 ;
        RECT  2.400 0.535 2.510 1.195 ;
        RECT  2.280 0.260 2.490 0.375 ;
        RECT  2.085 0.535 2.400 0.645 ;
        RECT  2.095 1.085 2.400 1.195 ;
        RECT  1.150 0.275 2.280 0.375 ;
        RECT  1.975 0.790 2.170 0.900 ;
        RECT  1.885 0.480 1.975 1.300 ;
        RECT  1.565 0.480 1.885 0.590 ;
        RECT  1.595 1.210 1.885 1.300 ;
        RECT  1.195 1.170 1.305 1.280 ;
        RECT  1.195 0.520 1.300 0.630 ;
        RECT  1.105 0.520 1.195 1.280 ;
        RECT  1.050 0.275 1.150 0.410 ;
        RECT  0.830 0.310 1.050 0.410 ;
        RECT  0.880 1.110 0.995 1.500 ;
        RECT  0.740 0.500 0.850 0.965 ;
        RECT  0.350 0.500 0.740 0.590 ;
        RECT  0.260 0.500 0.350 1.320 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.230 0.260 1.320 ;
        RECT  0.075 0.300 0.185 0.590 ;
        RECT  0.075 1.230 0.185 1.495 ;
    END
END DFXD2

MACRO DFXD4
    CLASS CORE ;
    FOREIGN DFXD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.275 7.265 0.675 ;
        RECT  7.250 1.040 7.265 1.470 ;
        RECT  7.155 0.275 7.250 1.470 ;
        RECT  6.950 0.505 7.155 1.210 ;
        RECT  6.765 0.505 6.950 0.675 ;
        RECT  6.765 1.040 6.950 1.210 ;
        RECT  6.655 0.275 6.765 0.675 ;
        RECT  6.655 1.040 6.765 1.470 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.545 6.295 0.655 ;
        RECT  6.135 1.040 6.245 1.470 ;
        RECT  6.050 1.040 6.135 1.140 ;
        RECT  5.750 0.545 6.050 1.140 ;
        RECT  5.565 0.545 5.750 0.655 ;
        RECT  5.725 1.040 5.750 1.140 ;
        RECT  5.615 1.040 5.725 1.470 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.315 0.750 1.450 0.920 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.590 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.760 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.525 -0.165 7.600 0.165 ;
        RECT  7.415 -0.165 7.525 0.695 ;
        RECT  3.265 -0.165 7.415 0.165 ;
        RECT  3.095 -0.165 3.265 0.295 ;
        RECT  0.480 -0.165 3.095 0.165 ;
        RECT  0.305 -0.165 0.480 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.525 1.635 7.600 1.965 ;
        RECT  7.415 1.040 7.525 1.965 ;
        RECT  6.505 1.635 7.415 1.965 ;
        RECT  6.395 1.040 6.505 1.965 ;
        RECT  5.985 1.635 6.395 1.965 ;
        RECT  5.875 1.260 5.985 1.965 ;
        RECT  5.465 1.635 5.875 1.965 ;
        RECT  5.355 1.040 5.465 1.965 ;
        RECT  3.200 1.635 5.355 1.965 ;
        RECT  3.200 1.195 3.320 1.305 ;
        RECT  3.085 1.195 3.200 1.965 ;
        RECT  0.500 1.635 3.085 1.965 ;
        RECT  0.330 1.415 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.765 0.505 6.850 0.675 ;
        RECT  6.765 1.040 6.850 1.210 ;
        RECT  6.655 0.275 6.765 0.675 ;
        RECT  6.655 1.040 6.765 1.470 ;
        RECT  6.150 0.545 6.295 0.655 ;
        RECT  6.150 1.040 6.245 1.470 ;
        RECT  5.565 0.545 5.650 0.655 ;
        RECT  5.615 1.040 5.650 1.470 ;
        RECT  6.545 0.780 6.720 0.890 ;
        RECT  6.435 0.345 6.545 0.890 ;
        RECT  4.200 0.345 6.435 0.455 ;
        RECT  5.265 0.780 5.600 0.890 ;
        RECT  5.205 0.545 5.265 1.140 ;
        RECT  5.170 0.545 5.205 1.470 ;
        RECT  4.470 0.545 5.170 0.655 ;
        RECT  5.095 1.040 5.170 1.470 ;
        RECT  4.895 0.750 5.005 1.525 ;
        RECT  3.810 1.435 4.895 1.525 ;
        RECT  4.230 1.085 4.770 1.195 ;
        RECT  4.360 0.545 4.470 0.940 ;
        RECT  4.200 1.085 4.230 1.275 ;
        RECT  4.100 0.345 4.200 1.275 ;
        RECT  4.000 0.275 4.010 1.030 ;
        RECT  3.910 0.275 4.000 1.245 ;
        RECT  3.570 0.275 3.910 0.365 ;
        RECT  3.900 0.930 3.910 1.245 ;
        RECT  3.810 0.455 3.820 0.820 ;
        RECT  3.710 0.455 3.810 1.525 ;
        RECT  3.700 0.710 3.710 1.525 ;
        RECT  3.480 0.275 3.570 0.475 ;
        RECT  3.455 0.565 3.555 1.255 ;
        RECT  2.935 0.385 3.480 0.475 ;
        RECT  3.105 0.565 3.455 0.665 ;
        RECT  3.255 0.765 3.365 1.105 ;
        RECT  2.765 1.015 3.255 1.105 ;
        RECT  2.995 0.565 3.105 0.925 ;
        RECT  2.825 0.275 2.935 0.475 ;
        RECT  2.715 1.015 2.765 1.340 ;
        RECT  2.655 0.415 2.715 1.340 ;
        RECT  2.615 0.415 2.655 1.105 ;
        RECT  0.995 1.390 2.520 1.500 ;
        RECT  2.400 0.535 2.510 1.195 ;
        RECT  1.150 0.275 2.495 0.375 ;
        RECT  2.085 0.535 2.400 0.645 ;
        RECT  2.095 1.085 2.400 1.195 ;
        RECT  1.975 0.790 2.170 0.900 ;
        RECT  1.885 0.480 1.975 1.300 ;
        RECT  1.565 0.480 1.885 0.590 ;
        RECT  1.595 1.210 1.885 1.300 ;
        RECT  1.195 1.170 1.305 1.280 ;
        RECT  1.195 0.520 1.300 0.630 ;
        RECT  1.105 0.520 1.195 1.280 ;
        RECT  1.050 0.275 1.150 0.410 ;
        RECT  0.830 0.310 1.050 0.410 ;
        RECT  0.880 1.110 0.995 1.500 ;
        RECT  0.740 0.500 0.850 0.965 ;
        RECT  0.350 0.500 0.740 0.590 ;
        RECT  0.260 0.500 0.350 1.320 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.230 0.260 1.320 ;
        RECT  0.075 0.300 0.185 0.590 ;
        RECT  0.075 1.230 0.185 1.495 ;
    END
END DFXD4

MACRO DFXQD1
    CLASS CORE ;
    FOREIGN DFXQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.275 4.950 1.490 ;
        RECT  4.825 0.275 4.850 0.660 ;
        RECT  4.815 1.020 4.850 1.490 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.550 1.090 ;
        RECT  1.315 0.750 1.450 0.920 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.590 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.710 1.765 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.480 -0.165 5.000 0.165 ;
        RECT  0.305 -0.165 0.480 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.195 1.635 5.000 1.965 ;
        RECT  3.020 1.355 3.195 1.965 ;
        RECT  0.475 1.635 3.020 1.965 ;
        RECT  0.305 1.415 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.670 0.750 4.760 0.920 ;
        RECT  4.570 0.525 4.670 1.420 ;
        RECT  4.390 0.525 4.570 0.615 ;
        RECT  4.260 1.310 4.570 1.420 ;
        RECT  4.305 0.780 4.460 0.890 ;
        RECT  4.280 0.275 4.390 0.615 ;
        RECT  4.215 0.780 4.305 1.160 ;
        RECT  4.070 0.525 4.280 0.615 ;
        RECT  4.125 1.070 4.215 1.160 ;
        RECT  4.035 1.070 4.125 1.495 ;
        RECT  3.980 0.525 4.070 0.960 ;
        RECT  3.655 1.395 4.035 1.495 ;
        RECT  3.840 0.275 3.880 0.950 ;
        RECT  3.790 0.275 3.840 1.285 ;
        RECT  3.575 0.275 3.790 0.365 ;
        RECT  3.750 0.835 3.790 1.285 ;
        RECT  3.655 0.465 3.700 0.660 ;
        RECT  3.565 0.465 3.655 1.495 ;
        RECT  3.365 0.255 3.575 0.365 ;
        RECT  3.545 1.395 3.565 1.495 ;
        RECT  3.370 0.475 3.475 1.245 ;
        RECT  3.250 0.475 3.370 0.585 ;
        RECT  3.040 1.135 3.370 1.245 ;
        RECT  2.865 0.275 3.365 0.365 ;
        RECT  3.175 0.700 3.280 1.005 ;
        RECT  2.700 0.700 3.175 0.790 ;
        RECT  2.925 0.900 3.040 1.245 ;
        RECT  2.665 0.255 2.865 0.365 ;
        RECT  2.690 0.500 2.700 0.790 ;
        RECT  2.570 0.500 2.690 1.330 ;
        RECT  2.250 0.275 2.470 0.385 ;
        RECT  2.320 0.535 2.450 1.195 ;
        RECT  0.930 1.420 2.440 1.525 ;
        RECT  2.060 0.535 2.320 0.670 ;
        RECT  2.060 1.065 2.320 1.195 ;
        RECT  1.040 0.275 2.250 0.370 ;
        RECT  1.950 0.770 2.105 0.900 ;
        RECT  1.860 0.500 1.950 1.290 ;
        RECT  1.580 0.500 1.860 0.600 ;
        RECT  1.555 1.200 1.860 1.290 ;
        RECT  1.130 0.520 1.300 0.630 ;
        RECT  1.130 1.170 1.250 1.280 ;
        RECT  1.040 0.520 1.130 1.280 ;
        RECT  0.830 0.275 1.040 0.410 ;
        RECT  0.820 1.110 0.930 1.525 ;
        RECT  0.715 0.500 0.830 0.965 ;
        RECT  0.350 0.500 0.715 0.590 ;
        RECT  0.260 0.500 0.350 1.320 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.230 0.260 1.320 ;
        RECT  0.075 0.300 0.185 0.590 ;
        RECT  0.075 1.230 0.185 1.495 ;
    END
END DFXQD1

MACRO DFXQD2
    CLASS CORE ;
    FOREIGN DFXQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.575 5.350 1.140 ;
        RECT  5.050 0.575 5.250 0.690 ;
        RECT  5.050 1.040 5.250 1.140 ;
        RECT  4.920 0.275 5.050 0.690 ;
        RECT  4.920 1.040 5.050 1.490 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.550 1.090 ;
        RECT  1.315 0.750 1.450 0.920 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.590 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.710 1.765 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.300 -0.165 5.400 0.165 ;
        RECT  5.190 -0.165 5.300 0.485 ;
        RECT  4.780 -0.165 5.190 0.165 ;
        RECT  4.670 -0.165 4.780 0.465 ;
        RECT  4.240 -0.165 4.670 0.165 ;
        RECT  4.110 -0.165 4.240 0.445 ;
        RECT  0.480 -0.165 4.110 0.165 ;
        RECT  0.305 -0.165 0.480 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.300 1.635 5.400 1.965 ;
        RECT  5.190 1.260 5.300 1.965 ;
        RECT  4.780 1.635 5.190 1.965 ;
        RECT  4.670 1.260 4.780 1.965 ;
        RECT  4.240 1.635 4.670 1.965 ;
        RECT  4.110 1.295 4.240 1.965 ;
        RECT  3.195 1.635 4.110 1.965 ;
        RECT  3.020 1.355 3.195 1.965 ;
        RECT  0.475 1.635 3.020 1.965 ;
        RECT  0.305 1.415 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.780 0.780 5.100 0.890 ;
        RECT  4.680 0.565 4.780 1.140 ;
        RECT  4.520 0.565 4.680 0.675 ;
        RECT  4.520 1.040 4.680 1.140 ;
        RECT  4.280 0.780 4.570 0.890 ;
        RECT  4.410 0.275 4.520 0.675 ;
        RECT  4.410 1.040 4.520 1.470 ;
        RECT  4.070 0.565 4.410 0.675 ;
        RECT  4.190 0.780 4.280 1.185 ;
        RECT  4.020 1.095 4.190 1.185 ;
        RECT  3.980 0.565 4.070 0.960 ;
        RECT  3.930 1.095 4.020 1.495 ;
        RECT  3.655 1.395 3.930 1.495 ;
        RECT  3.840 0.275 3.880 0.950 ;
        RECT  3.790 0.275 3.840 1.285 ;
        RECT  3.575 0.275 3.790 0.365 ;
        RECT  3.750 0.835 3.790 1.285 ;
        RECT  3.655 0.465 3.700 0.660 ;
        RECT  3.565 0.465 3.655 1.495 ;
        RECT  3.365 0.255 3.575 0.365 ;
        RECT  3.545 1.395 3.565 1.495 ;
        RECT  3.370 0.475 3.475 1.245 ;
        RECT  3.250 0.475 3.370 0.585 ;
        RECT  3.040 1.135 3.370 1.245 ;
        RECT  2.865 0.275 3.365 0.365 ;
        RECT  3.175 0.700 3.280 1.005 ;
        RECT  2.700 0.700 3.175 0.790 ;
        RECT  2.925 0.900 3.040 1.245 ;
        RECT  2.665 0.255 2.865 0.365 ;
        RECT  2.690 0.500 2.700 0.790 ;
        RECT  2.570 0.500 2.690 1.330 ;
        RECT  2.250 0.275 2.460 0.385 ;
        RECT  2.320 0.535 2.450 1.195 ;
        RECT  0.930 1.420 2.440 1.525 ;
        RECT  2.060 0.535 2.320 0.670 ;
        RECT  2.060 1.065 2.320 1.195 ;
        RECT  1.040 0.275 2.250 0.370 ;
        RECT  1.950 0.770 2.105 0.900 ;
        RECT  1.860 0.500 1.950 1.290 ;
        RECT  1.580 0.500 1.860 0.600 ;
        RECT  1.555 1.200 1.860 1.290 ;
        RECT  1.130 0.520 1.300 0.630 ;
        RECT  1.130 1.170 1.250 1.280 ;
        RECT  1.040 0.520 1.130 1.280 ;
        RECT  0.830 0.275 1.040 0.410 ;
        RECT  0.820 1.110 0.930 1.525 ;
        RECT  0.715 0.500 0.830 0.965 ;
        RECT  0.350 0.500 0.715 0.590 ;
        RECT  0.260 0.500 0.350 1.320 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.230 0.260 1.320 ;
        RECT  0.075 0.300 0.185 0.590 ;
        RECT  0.075 1.230 0.185 1.495 ;
    END
END DFXQD2

MACRO DFXQD4
    CLASS CORE ;
    FOREIGN DFXQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.275 5.675 0.675 ;
        RECT  5.650 1.040 5.675 1.470 ;
        RECT  5.555 0.275 5.650 1.470 ;
        RECT  5.545 0.275 5.555 1.140 ;
        RECT  5.325 0.575 5.545 1.140 ;
        RECT  5.145 0.575 5.325 0.675 ;
        RECT  5.145 1.040 5.325 1.140 ;
        RECT  5.035 0.275 5.145 0.675 ;
        RECT  5.035 1.040 5.145 1.470 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.315 0.750 1.450 0.920 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0328 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.590 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.760 1.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.940 -0.165 6.000 0.165 ;
        RECT  5.805 -0.165 5.940 0.705 ;
        RECT  5.420 -0.165 5.805 0.165 ;
        RECT  5.285 -0.165 5.420 0.465 ;
        RECT  4.895 -0.165 5.285 0.165 ;
        RECT  4.765 -0.165 4.895 0.465 ;
        RECT  4.355 -0.165 4.765 0.165 ;
        RECT  4.230 -0.165 4.355 0.465 ;
        RECT  3.265 -0.165 4.230 0.165 ;
        RECT  3.095 -0.165 3.265 0.295 ;
        RECT  0.480 -0.165 3.095 0.165 ;
        RECT  0.305 -0.165 0.480 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.935 1.635 6.000 1.965 ;
        RECT  5.805 1.035 5.935 1.965 ;
        RECT  5.415 1.635 5.805 1.965 ;
        RECT  5.285 1.295 5.415 1.965 ;
        RECT  4.885 1.635 5.285 1.965 ;
        RECT  4.775 1.260 4.885 1.965 ;
        RECT  3.200 1.635 4.775 1.965 ;
        RECT  3.200 1.195 3.320 1.305 ;
        RECT  3.085 1.195 3.200 1.965 ;
        RECT  0.500 1.635 3.085 1.965 ;
        RECT  0.330 1.415 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.145 0.575 5.250 0.675 ;
        RECT  5.145 1.040 5.250 1.140 ;
        RECT  5.035 0.275 5.145 0.675 ;
        RECT  5.035 1.040 5.145 1.470 ;
        RECT  4.885 0.780 5.175 0.890 ;
        RECT  4.785 0.565 4.885 1.140 ;
        RECT  4.625 0.565 4.785 0.675 ;
        RECT  4.625 1.040 4.785 1.140 ;
        RECT  4.380 0.780 4.675 0.890 ;
        RECT  4.515 0.275 4.625 0.675 ;
        RECT  4.515 1.040 4.625 1.470 ;
        RECT  4.200 0.565 4.515 0.675 ;
        RECT  4.290 0.780 4.380 1.495 ;
        RECT  3.810 1.385 4.290 1.495 ;
        RECT  4.110 0.565 4.200 0.940 ;
        RECT  3.920 0.275 4.020 1.265 ;
        RECT  3.570 0.275 3.920 0.365 ;
        RECT  3.900 1.055 3.920 1.265 ;
        RECT  3.810 0.455 3.830 0.645 ;
        RECT  3.700 0.455 3.810 1.495 ;
        RECT  3.655 1.385 3.700 1.495 ;
        RECT  3.480 0.275 3.570 0.475 ;
        RECT  3.455 0.565 3.555 1.255 ;
        RECT  2.935 0.385 3.480 0.475 ;
        RECT  3.105 0.565 3.455 0.665 ;
        RECT  3.255 0.765 3.365 1.105 ;
        RECT  2.765 1.015 3.255 1.105 ;
        RECT  2.995 0.565 3.105 0.925 ;
        RECT  2.825 0.275 2.935 0.475 ;
        RECT  2.715 1.015 2.765 1.340 ;
        RECT  2.655 0.415 2.715 1.340 ;
        RECT  2.615 0.415 2.655 1.105 ;
        RECT  2.355 1.370 2.520 1.480 ;
        RECT  2.400 0.535 2.510 1.195 ;
        RECT  1.150 0.275 2.495 0.375 ;
        RECT  2.085 0.535 2.400 0.645 ;
        RECT  2.095 1.085 2.400 1.195 ;
        RECT  2.245 1.370 2.355 1.525 ;
        RECT  0.995 1.415 2.245 1.525 ;
        RECT  1.975 0.790 2.170 0.900 ;
        RECT  1.885 0.480 1.975 1.320 ;
        RECT  1.565 0.480 1.885 0.590 ;
        RECT  1.595 1.210 1.885 1.320 ;
        RECT  1.195 1.170 1.305 1.280 ;
        RECT  1.195 0.520 1.300 0.630 ;
        RECT  1.105 0.520 1.195 1.280 ;
        RECT  1.050 0.275 1.150 0.410 ;
        RECT  0.830 0.310 1.050 0.410 ;
        RECT  0.880 1.130 0.995 1.525 ;
        RECT  0.740 0.500 0.850 0.965 ;
        RECT  0.350 0.500 0.740 0.590 ;
        RECT  0.260 0.500 0.350 1.320 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.230 0.260 1.320 ;
        RECT  0.075 0.300 0.185 0.590 ;
        RECT  0.075 1.230 0.185 1.495 ;
    END
END DFXQD4

MACRO EDFCND1
    CLASS CORE ;
    FOREIGN EDFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.275 6.150 1.490 ;
        RECT  6.020 0.275 6.050 0.675 ;
        RECT  6.020 1.040 6.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.575 5.750 1.300 ;
        RECT  5.600 0.575 5.650 0.675 ;
        RECT  5.480 1.090 5.650 1.300 ;
        RECT  5.480 0.285 5.600 0.675 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0661 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.710 1.750 0.910 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0669 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.510 4.970 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.870 -0.165 6.200 0.165 ;
        RECT  5.740 -0.165 5.870 0.470 ;
        RECT  4.565 -0.165 5.740 0.165 ;
        RECT  4.395 -0.165 4.565 0.385 ;
        RECT  3.395 -0.165 4.395 0.165 ;
        RECT  3.285 -0.165 3.395 0.405 ;
        RECT  0.560 -0.165 3.285 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.635 6.200 1.965 ;
        RECT  3.245 1.445 3.415 1.965 ;
        RECT  0.475 1.635 3.245 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.930 0.755 5.945 0.925 ;
        RECT  5.840 0.755 5.930 1.515 ;
        RECT  4.490 1.425 5.840 1.515 ;
        RECT  5.375 0.765 5.435 0.935 ;
        RECT  5.275 0.285 5.375 1.305 ;
        RECT  5.240 0.285 5.275 0.675 ;
        RECT  4.690 1.200 5.275 1.305 ;
        RECT  5.150 0.765 5.185 0.935 ;
        RECT  5.060 0.315 5.150 0.935 ;
        RECT  4.745 0.315 5.060 0.415 ;
        RECT  4.655 0.315 4.745 0.585 ;
        RECT  4.580 0.875 4.690 1.305 ;
        RECT  4.490 0.675 4.670 0.765 ;
        RECT  4.040 0.495 4.655 0.585 ;
        RECT  4.380 0.675 4.490 1.515 ;
        RECT  4.150 0.675 4.380 0.765 ;
        RECT  3.605 1.425 4.380 1.515 ;
        RECT  4.075 0.865 4.185 1.315 ;
        RECT  4.040 0.865 4.075 0.975 ;
        RECT  3.940 0.495 4.040 0.975 ;
        RECT  3.575 0.305 3.965 0.405 ;
        RECT  3.815 1.085 3.920 1.315 ;
        RECT  3.795 1.085 3.815 1.175 ;
        RECT  3.680 0.495 3.795 1.175 ;
        RECT  3.665 0.905 3.680 1.175 ;
        RECT  2.900 0.905 3.665 0.995 ;
        RECT  3.505 1.265 3.605 1.515 ;
        RECT  2.700 0.705 3.590 0.815 ;
        RECT  3.485 0.305 3.575 0.585 ;
        RECT  3.155 1.265 3.505 1.355 ;
        RECT  3.065 0.495 3.485 0.585 ;
        RECT  2.945 1.085 3.455 1.175 ;
        RECT  3.065 1.265 3.155 1.525 ;
        RECT  2.975 0.280 3.065 0.585 ;
        RECT  2.600 1.435 3.065 1.525 ;
        RECT  2.675 0.280 2.975 0.390 ;
        RECT  2.775 1.085 2.945 1.310 ;
        RECT  2.665 0.495 2.700 0.815 ;
        RECT  2.575 0.495 2.665 1.140 ;
        RECT  2.510 1.255 2.600 1.525 ;
        RECT  2.475 1.030 2.575 1.140 ;
        RECT  1.340 1.255 2.510 1.345 ;
        RECT  1.035 0.275 2.465 0.385 ;
        RECT  1.085 1.435 2.400 1.525 ;
        RECT  2.220 0.510 2.330 1.145 ;
        RECT  2.025 0.510 2.220 0.645 ;
        RECT  2.030 1.025 2.220 1.145 ;
        RECT  1.930 0.785 2.105 0.905 ;
        RECT  1.840 0.490 1.930 1.145 ;
        RECT  1.530 0.490 1.840 0.600 ;
        RECT  1.500 1.030 1.840 1.145 ;
        RECT  1.230 0.915 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFCND1

MACRO EDFCND2
    CLASS CORE ;
    FOREIGN EDFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.655 0.595 6.750 1.150 ;
        RECT  6.605 0.595 6.655 0.695 ;
        RECT  6.625 1.040 6.655 1.150 ;
        RECT  6.450 1.040 6.625 1.490 ;
        RECT  6.450 0.275 6.605 0.695 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.015 0.285 6.150 1.300 ;
        RECT  5.970 0.285 6.015 0.675 ;
        RECT  5.970 1.045 6.015 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0661 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.710 1.750 0.910 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0995 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.510 4.970 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.880 -0.165 7.000 0.165 ;
        RECT  6.755 -0.165 6.880 0.485 ;
        RECT  6.360 -0.165 6.755 0.165 ;
        RECT  6.250 -0.165 6.360 0.675 ;
        RECT  5.825 -0.165 6.250 0.165 ;
        RECT  5.700 -0.165 5.825 0.675 ;
        RECT  4.565 -0.165 5.700 0.165 ;
        RECT  4.395 -0.165 4.565 0.355 ;
        RECT  3.395 -0.165 4.395 0.165 ;
        RECT  3.285 -0.165 3.395 0.405 ;
        RECT  0.560 -0.165 3.285 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.880 1.635 7.000 1.965 ;
        RECT  6.755 1.260 6.880 1.965 ;
        RECT  3.415 1.635 6.755 1.965 ;
        RECT  3.245 1.445 3.415 1.965 ;
        RECT  0.475 1.635 3.245 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.350 0.785 6.530 0.895 ;
        RECT  6.250 0.785 6.350 1.515 ;
        RECT  4.490 1.425 6.250 1.515 ;
        RECT  5.580 0.765 5.925 0.935 ;
        RECT  5.470 0.545 5.580 1.305 ;
        RECT  5.160 0.545 5.470 0.655 ;
        RECT  4.690 1.200 5.470 1.305 ;
        RECT  4.745 0.305 5.400 0.405 ;
        RECT  4.655 0.305 4.745 0.585 ;
        RECT  4.580 0.875 4.690 1.305 ;
        RECT  4.490 0.675 4.670 0.765 ;
        RECT  4.040 0.495 4.655 0.585 ;
        RECT  4.380 0.675 4.490 1.515 ;
        RECT  4.150 0.675 4.380 0.765 ;
        RECT  3.605 1.425 4.380 1.515 ;
        RECT  4.075 0.865 4.185 1.315 ;
        RECT  4.040 0.865 4.075 0.975 ;
        RECT  3.940 0.495 4.040 0.975 ;
        RECT  3.575 0.305 3.965 0.405 ;
        RECT  3.815 1.085 3.920 1.315 ;
        RECT  3.795 1.085 3.815 1.175 ;
        RECT  3.680 0.495 3.795 1.175 ;
        RECT  3.665 0.905 3.680 1.175 ;
        RECT  2.900 0.905 3.665 0.995 ;
        RECT  3.505 1.265 3.605 1.515 ;
        RECT  2.700 0.705 3.590 0.815 ;
        RECT  3.485 0.305 3.575 0.585 ;
        RECT  3.155 1.265 3.505 1.355 ;
        RECT  3.065 0.495 3.485 0.585 ;
        RECT  2.945 1.085 3.455 1.175 ;
        RECT  3.065 1.265 3.155 1.525 ;
        RECT  2.975 0.280 3.065 0.585 ;
        RECT  2.600 1.435 3.065 1.525 ;
        RECT  2.675 0.280 2.975 0.390 ;
        RECT  2.775 1.085 2.945 1.310 ;
        RECT  2.665 0.495 2.700 0.815 ;
        RECT  2.575 0.495 2.665 1.140 ;
        RECT  2.510 1.255 2.600 1.525 ;
        RECT  2.475 1.030 2.575 1.140 ;
        RECT  1.340 1.255 2.510 1.345 ;
        RECT  1.035 0.275 2.465 0.385 ;
        RECT  1.085 1.435 2.400 1.525 ;
        RECT  2.220 0.510 2.330 1.145 ;
        RECT  2.025 0.510 2.220 0.645 ;
        RECT  2.030 1.025 2.220 1.145 ;
        RECT  1.930 0.785 2.105 0.905 ;
        RECT  1.840 0.490 1.930 1.145 ;
        RECT  1.530 0.490 1.840 0.600 ;
        RECT  1.500 1.030 1.840 1.145 ;
        RECT  1.230 0.915 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFCND2

MACRO EDFCND4
    CLASS CORE ;
    FOREIGN EDFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 0.315 8.095 0.645 ;
        RECT  7.850 1.060 8.095 1.430 ;
        RECT  7.560 0.315 7.850 1.430 ;
        RECT  7.415 0.315 7.560 0.645 ;
        RECT  7.415 1.060 7.560 1.430 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.475 7.085 0.675 ;
        RECT  6.850 1.040 7.085 1.290 ;
        RECT  6.550 0.475 6.850 1.290 ;
        RECT  6.415 0.475 6.550 0.675 ;
        RECT  6.415 1.040 6.550 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0643 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.910 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0991 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.845 0.510 4.965 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.330 -0.165 8.400 0.165 ;
        RECT  8.210 -0.165 8.330 0.685 ;
        RECT  5.785 -0.165 8.210 0.165 ;
        RECT  5.675 -0.165 5.785 0.645 ;
        RECT  4.560 -0.165 5.675 0.165 ;
        RECT  4.390 -0.165 4.560 0.355 ;
        RECT  3.390 -0.165 4.390 0.165 ;
        RECT  3.280 -0.165 3.390 0.405 ;
        RECT  0.560 -0.165 3.280 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.330 1.635 8.400 1.965 ;
        RECT  8.210 1.030 8.330 1.965 ;
        RECT  3.410 1.635 8.210 1.965 ;
        RECT  3.240 1.445 3.410 1.965 ;
        RECT  0.475 1.635 3.240 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.950 0.315 8.095 0.645 ;
        RECT  7.950 1.060 8.095 1.430 ;
        RECT  7.415 0.315 7.450 0.645 ;
        RECT  7.415 1.060 7.450 1.430 ;
        RECT  6.960 0.475 7.085 0.675 ;
        RECT  6.960 1.040 7.085 1.290 ;
        RECT  6.415 0.475 6.460 0.675 ;
        RECT  6.415 1.040 6.460 1.290 ;
        RECT  7.315 0.765 7.450 0.935 ;
        RECT  7.310 0.765 7.315 1.515 ;
        RECT  7.195 0.275 7.310 1.515 ;
        RECT  6.065 0.275 7.195 0.365 ;
        RECT  6.060 1.410 7.195 1.515 ;
        RECT  5.575 0.785 6.440 0.915 ;
        RECT  5.935 0.275 6.065 0.655 ;
        RECT  5.940 1.060 6.060 1.515 ;
        RECT  4.485 1.410 5.940 1.515 ;
        RECT  5.465 0.545 5.575 1.305 ;
        RECT  5.155 0.545 5.465 0.655 ;
        RECT  4.685 1.200 5.465 1.305 ;
        RECT  4.740 0.315 5.395 0.405 ;
        RECT  4.650 0.315 4.740 0.585 ;
        RECT  4.575 0.875 4.685 1.305 ;
        RECT  4.485 0.675 4.665 0.765 ;
        RECT  4.035 0.495 4.650 0.585 ;
        RECT  4.375 0.675 4.485 1.515 ;
        RECT  4.145 0.675 4.375 0.765 ;
        RECT  3.600 1.425 4.375 1.515 ;
        RECT  4.070 0.865 4.180 1.315 ;
        RECT  4.035 0.865 4.070 0.975 ;
        RECT  3.935 0.495 4.035 0.975 ;
        RECT  3.570 0.305 3.960 0.405 ;
        RECT  3.810 1.085 3.915 1.315 ;
        RECT  3.790 1.085 3.810 1.175 ;
        RECT  3.675 0.495 3.790 1.175 ;
        RECT  3.660 0.905 3.675 1.175 ;
        RECT  2.895 0.905 3.660 0.995 ;
        RECT  3.500 1.265 3.600 1.515 ;
        RECT  2.695 0.705 3.585 0.815 ;
        RECT  3.480 0.305 3.570 0.585 ;
        RECT  3.150 1.265 3.500 1.355 ;
        RECT  3.060 0.495 3.480 0.585 ;
        RECT  2.940 1.085 3.450 1.175 ;
        RECT  3.060 1.265 3.150 1.525 ;
        RECT  2.970 0.280 3.060 0.585 ;
        RECT  2.595 1.435 3.060 1.525 ;
        RECT  2.670 0.280 2.970 0.390 ;
        RECT  2.770 1.085 2.940 1.310 ;
        RECT  2.660 0.495 2.695 0.815 ;
        RECT  2.570 0.495 2.660 1.140 ;
        RECT  2.505 1.255 2.595 1.525 ;
        RECT  2.470 1.030 2.570 1.140 ;
        RECT  1.340 1.255 2.505 1.345 ;
        RECT  1.035 0.275 2.460 0.385 ;
        RECT  1.085 1.435 2.395 1.525 ;
        RECT  2.215 0.510 2.325 1.145 ;
        RECT  2.020 0.510 2.215 0.645 ;
        RECT  2.020 1.025 2.215 1.145 ;
        RECT  1.930 0.785 2.090 0.905 ;
        RECT  1.840 0.490 1.930 1.145 ;
        RECT  1.515 0.490 1.840 0.600 ;
        RECT  1.485 1.030 1.840 1.145 ;
        RECT  1.235 0.900 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFCND4

MACRO EDFCNQD1
    CLASS CORE ;
    FOREIGN EDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.665 0.585 5.755 1.150 ;
        RECT  5.645 0.285 5.665 1.470 ;
        RECT  5.555 0.285 5.645 0.695 ;
        RECT  5.555 1.040 5.645 1.470 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0689 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.355 1.120 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.750 0.600 0.920 ;
        RECT  0.445 0.510 0.555 0.920 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.690 1.620 0.890 ;
        RECT  1.355 0.690 1.450 0.800 ;
        RECT  1.245 0.480 1.355 0.800 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0575 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.045 0.480 5.155 1.030 ;
        RECT  4.910 0.850 5.045 1.030 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.925 -0.165 6.000 0.165 ;
        RECT  5.815 -0.165 5.925 0.475 ;
        RECT  4.745 -0.165 5.815 0.165 ;
        RECT  4.575 -0.165 4.745 0.355 ;
        RECT  3.400 -0.165 4.575 0.165 ;
        RECT  3.290 -0.165 3.400 0.405 ;
        RECT  0.485 -0.165 3.290 0.165 ;
        RECT  0.315 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.925 1.635 6.000 1.965 ;
        RECT  5.815 1.260 5.925 1.965 ;
        RECT  5.375 1.635 5.815 1.965 ;
        RECT  5.265 1.335 5.375 1.965 ;
        RECT  3.680 1.635 5.265 1.965 ;
        RECT  3.510 1.445 3.680 1.965 ;
        RECT  0.585 1.635 3.510 1.965 ;
        RECT  0.475 1.395 0.585 1.965 ;
        RECT  0.285 1.395 0.475 1.505 ;
        RECT  0.000 1.635 0.475 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.380 0.785 5.535 0.890 ;
        RECT  5.265 0.460 5.380 1.245 ;
        RECT  4.935 0.275 5.345 0.365 ;
        RECT  5.115 1.130 5.265 1.245 ;
        RECT  5.005 1.130 5.115 1.515 ;
        RECT  4.800 1.130 5.005 1.245 ;
        RECT  4.845 0.275 4.935 0.535 ;
        RECT  4.310 0.445 4.845 0.535 ;
        RECT  4.690 0.900 4.800 1.245 ;
        RECT  4.515 0.635 4.715 0.745 ;
        RECT  4.605 0.900 4.690 1.010 ;
        RECT  4.515 1.115 4.595 1.515 ;
        RECT  4.425 0.635 4.515 1.515 ;
        RECT  4.215 0.685 4.425 0.775 ;
        RECT  3.870 1.425 4.425 1.515 ;
        RECT  4.225 0.865 4.335 1.305 ;
        RECT  4.200 0.445 4.310 0.595 ;
        RECT  4.105 0.865 4.225 0.975 ;
        RECT  4.105 0.505 4.200 0.595 ;
        RECT  3.990 0.505 4.105 0.975 ;
        RECT  3.965 1.065 4.075 1.315 ;
        RECT  3.580 0.305 4.010 0.415 ;
        RECT  3.890 1.065 3.965 1.155 ;
        RECT  3.800 0.505 3.890 1.155 ;
        RECT  3.770 1.265 3.870 1.515 ;
        RECT  3.670 0.505 3.800 0.615 ;
        RECT  3.040 0.905 3.800 0.995 ;
        RECT  3.420 1.265 3.770 1.355 ;
        RECT  2.770 0.705 3.700 0.815 ;
        RECT  3.240 1.085 3.640 1.175 ;
        RECT  3.490 0.305 3.580 0.585 ;
        RECT  3.065 0.495 3.490 0.585 ;
        RECT  3.330 1.265 3.420 1.525 ;
        RECT  2.785 1.435 3.330 1.525 ;
        RECT  3.130 1.085 3.240 1.310 ;
        RECT  2.940 1.200 3.130 1.310 ;
        RECT  2.975 0.280 3.065 0.585 ;
        RECT  2.870 0.905 3.040 1.050 ;
        RECT  2.690 0.280 2.975 0.390 ;
        RECT  2.695 1.255 2.785 1.525 ;
        RECT  2.760 0.495 2.770 0.815 ;
        RECT  2.650 0.495 2.760 1.155 ;
        RECT  1.360 1.255 2.695 1.345 ;
        RECT  2.580 0.495 2.650 0.645 ;
        RECT  1.070 1.435 2.525 1.525 ;
        RECT  2.210 0.255 2.420 0.365 ;
        RECT  2.255 0.545 2.365 1.155 ;
        RECT  2.070 0.545 2.255 0.655 ;
        RECT  2.100 1.045 2.255 1.155 ;
        RECT  1.030 0.275 2.210 0.365 ;
        RECT  1.815 0.780 2.085 0.890 ;
        RECT  1.710 0.480 1.815 1.145 ;
        RECT  1.560 0.480 1.710 0.580 ;
        RECT  1.615 1.035 1.710 1.145 ;
        RECT  1.270 0.915 1.360 1.345 ;
        RECT  1.015 0.685 1.125 1.305 ;
        RECT  0.865 1.395 1.070 1.525 ;
        RECT  0.920 0.275 1.030 0.495 ;
        RECT  0.190 1.215 1.015 1.305 ;
        RECT  0.710 0.465 0.820 1.125 ;
        RECT  0.645 0.465 0.710 0.640 ;
        RECT  0.570 1.025 0.710 1.125 ;
        RECT  0.135 0.305 0.225 0.420 ;
        RECT  0.135 1.215 0.190 1.495 ;
        RECT  0.070 0.305 0.135 1.495 ;
        RECT  0.045 0.305 0.070 1.305 ;
    END
END EDFCNQD1

MACRO EDFCNQD2
    CLASS CORE ;
    FOREIGN EDFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.585 6.350 1.150 ;
        RECT  6.170 0.585 6.250 0.695 ;
        RECT  6.165 1.040 6.250 1.150 ;
        RECT  6.050 0.275 6.170 0.695 ;
        RECT  6.050 1.040 6.165 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0689 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.355 1.120 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.750 0.600 0.920 ;
        RECT  0.445 0.510 0.555 0.920 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.690 1.620 0.890 ;
        RECT  1.355 0.690 1.450 0.800 ;
        RECT  1.245 0.480 1.355 0.800 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0982 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.045 0.510 5.155 1.000 ;
        RECT  4.890 0.890 5.045 1.000 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.425 -0.165 6.600 0.165 ;
        RECT  6.315 -0.165 6.425 0.475 ;
        RECT  5.905 -0.165 6.315 0.165 ;
        RECT  5.795 -0.165 5.905 0.675 ;
        RECT  4.640 -0.165 5.795 0.165 ;
        RECT  4.470 -0.165 4.640 0.355 ;
        RECT  3.400 -0.165 4.470 0.165 ;
        RECT  3.290 -0.165 3.400 0.405 ;
        RECT  0.485 -0.165 3.290 0.165 ;
        RECT  0.315 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.425 1.635 6.600 1.965 ;
        RECT  6.315 1.260 6.425 1.965 ;
        RECT  5.905 1.635 6.315 1.965 ;
        RECT  5.795 1.040 5.905 1.965 ;
        RECT  5.385 1.635 5.795 1.965 ;
        RECT  5.275 1.330 5.385 1.965 ;
        RECT  3.680 1.635 5.275 1.965 ;
        RECT  3.510 1.445 3.680 1.965 ;
        RECT  0.585 1.635 3.510 1.965 ;
        RECT  0.475 1.395 0.585 1.965 ;
        RECT  0.285 1.395 0.475 1.505 ;
        RECT  0.000 1.635 0.475 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.645 0.785 6.140 0.895 ;
        RECT  5.535 0.785 5.645 1.515 ;
        RECT  5.385 0.785 5.535 0.895 ;
        RECT  5.125 1.130 5.535 1.240 ;
        RECT  4.935 0.315 5.415 0.420 ;
        RECT  5.275 0.510 5.385 0.895 ;
        RECT  5.015 1.130 5.125 1.515 ;
        RECT  4.800 1.130 5.015 1.240 ;
        RECT  4.845 0.315 4.935 0.535 ;
        RECT  4.310 0.445 4.845 0.535 ;
        RECT  4.690 0.900 4.800 1.240 ;
        RECT  4.515 0.625 4.715 0.735 ;
        RECT  4.605 0.900 4.690 1.010 ;
        RECT  4.515 1.115 4.595 1.515 ;
        RECT  4.425 0.625 4.515 1.515 ;
        RECT  4.215 0.685 4.425 0.775 ;
        RECT  3.870 1.425 4.425 1.515 ;
        RECT  4.225 0.865 4.335 1.305 ;
        RECT  4.200 0.445 4.310 0.595 ;
        RECT  4.105 0.865 4.225 0.975 ;
        RECT  4.105 0.505 4.200 0.595 ;
        RECT  3.990 0.505 4.105 0.975 ;
        RECT  3.965 1.065 4.075 1.315 ;
        RECT  3.580 0.305 4.010 0.415 ;
        RECT  3.890 1.065 3.965 1.155 ;
        RECT  3.800 0.505 3.890 1.155 ;
        RECT  3.770 1.265 3.870 1.515 ;
        RECT  3.670 0.505 3.800 0.615 ;
        RECT  3.040 0.905 3.800 0.995 ;
        RECT  3.420 1.265 3.770 1.355 ;
        RECT  2.770 0.705 3.700 0.815 ;
        RECT  3.240 1.085 3.640 1.175 ;
        RECT  3.490 0.305 3.580 0.585 ;
        RECT  3.065 0.495 3.490 0.585 ;
        RECT  3.330 1.265 3.420 1.525 ;
        RECT  2.785 1.435 3.330 1.525 ;
        RECT  3.130 1.085 3.240 1.310 ;
        RECT  2.940 1.200 3.130 1.310 ;
        RECT  2.975 0.280 3.065 0.585 ;
        RECT  2.870 0.905 3.040 1.050 ;
        RECT  2.690 0.280 2.975 0.390 ;
        RECT  2.695 1.255 2.785 1.525 ;
        RECT  2.760 0.495 2.770 0.815 ;
        RECT  2.650 0.495 2.760 1.155 ;
        RECT  1.360 1.255 2.695 1.345 ;
        RECT  2.580 0.495 2.650 0.645 ;
        RECT  1.070 1.435 2.525 1.525 ;
        RECT  2.210 0.255 2.420 0.365 ;
        RECT  2.255 0.545 2.365 1.155 ;
        RECT  2.035 0.545 2.255 0.655 ;
        RECT  2.110 1.045 2.255 1.155 ;
        RECT  1.030 0.275 2.210 0.365 ;
        RECT  1.815 0.780 2.085 0.890 ;
        RECT  1.710 0.480 1.815 1.145 ;
        RECT  1.560 0.480 1.710 0.580 ;
        RECT  1.615 1.035 1.710 1.145 ;
        RECT  1.270 0.915 1.360 1.345 ;
        RECT  1.015 0.685 1.125 1.305 ;
        RECT  0.865 1.395 1.070 1.525 ;
        RECT  0.920 0.275 1.030 0.495 ;
        RECT  0.190 1.215 1.015 1.305 ;
        RECT  0.710 0.465 0.820 1.125 ;
        RECT  0.645 0.465 0.710 0.640 ;
        RECT  0.570 1.025 0.710 1.125 ;
        RECT  0.135 0.305 0.225 0.420 ;
        RECT  0.135 1.215 0.190 1.495 ;
        RECT  0.070 0.305 0.135 1.495 ;
        RECT  0.045 0.305 0.070 1.305 ;
    END
END EDFCNQD2

MACRO EDFCNQD4
    CLASS CORE ;
    FOREIGN EDFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.495 6.645 0.690 ;
        RECT  6.450 1.040 6.645 1.290 ;
        RECT  6.150 0.495 6.450 1.290 ;
        RECT  5.955 0.495 6.150 0.690 ;
        RECT  5.955 1.040 6.150 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.800 1.695 0.910 ;
        RECT  1.450 0.690 1.550 0.910 ;
        RECT  1.370 0.690 1.450 0.790 ;
        RECT  1.245 0.510 1.370 0.790 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0996 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.845 0.510 4.965 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.885 -0.165 7.000 0.165 ;
        RECT  6.760 -0.165 6.885 0.705 ;
        RECT  6.385 -0.165 6.760 0.165 ;
        RECT  6.215 -0.165 6.385 0.405 ;
        RECT  5.845 -0.165 6.215 0.165 ;
        RECT  5.715 -0.165 5.845 0.645 ;
        RECT  4.560 -0.165 5.715 0.165 ;
        RECT  4.390 -0.165 4.560 0.385 ;
        RECT  3.390 -0.165 4.390 0.165 ;
        RECT  3.280 -0.165 3.390 0.405 ;
        RECT  0.560 -0.165 3.280 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.885 1.635 7.000 1.965 ;
        RECT  6.755 1.015 6.885 1.965 ;
        RECT  6.385 1.635 6.755 1.965 ;
        RECT  6.215 1.395 6.385 1.965 ;
        RECT  5.845 1.635 6.215 1.965 ;
        RECT  5.715 1.015 5.845 1.965 ;
        RECT  5.345 1.635 5.715 1.965 ;
        RECT  5.175 1.395 5.345 1.965 ;
        RECT  4.815 1.635 5.175 1.965 ;
        RECT  4.645 1.395 4.815 1.965 ;
        RECT  3.410 1.635 4.645 1.965 ;
        RECT  3.240 1.445 3.410 1.965 ;
        RECT  0.475 1.635 3.240 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.550 0.495 6.645 0.690 ;
        RECT  6.550 1.040 6.645 1.290 ;
        RECT  5.955 0.495 6.050 0.690 ;
        RECT  5.955 1.040 6.050 1.290 ;
        RECT  5.575 0.785 5.990 0.915 ;
        RECT  5.465 0.545 5.575 1.480 ;
        RECT  5.155 0.545 5.465 0.655 ;
        RECT  4.720 1.200 5.465 1.305 ;
        RECT  4.740 0.315 5.395 0.405 ;
        RECT  4.650 0.315 4.740 0.585 ;
        RECT  4.595 0.875 4.720 1.305 ;
        RECT  4.485 0.675 4.665 0.765 ;
        RECT  4.035 0.495 4.650 0.585 ;
        RECT  4.375 0.675 4.485 1.515 ;
        RECT  4.145 0.675 4.375 0.765 ;
        RECT  3.600 1.425 4.375 1.515 ;
        RECT  4.070 0.865 4.180 1.315 ;
        RECT  4.035 0.865 4.070 0.975 ;
        RECT  3.935 0.495 4.035 0.975 ;
        RECT  3.570 0.305 3.960 0.405 ;
        RECT  3.810 1.085 3.915 1.315 ;
        RECT  3.790 1.085 3.810 1.175 ;
        RECT  3.675 0.495 3.790 1.175 ;
        RECT  3.660 0.905 3.675 1.175 ;
        RECT  2.895 0.905 3.660 0.995 ;
        RECT  3.500 1.265 3.600 1.515 ;
        RECT  2.695 0.705 3.585 0.815 ;
        RECT  3.480 0.305 3.570 0.585 ;
        RECT  3.150 1.265 3.500 1.355 ;
        RECT  3.060 0.495 3.480 0.585 ;
        RECT  2.940 1.085 3.450 1.175 ;
        RECT  3.060 1.265 3.150 1.525 ;
        RECT  2.970 0.280 3.060 0.585 ;
        RECT  2.595 1.435 3.060 1.525 ;
        RECT  2.670 0.280 2.970 0.390 ;
        RECT  2.770 1.085 2.940 1.310 ;
        RECT  2.660 0.495 2.695 0.815 ;
        RECT  2.570 0.495 2.660 1.140 ;
        RECT  2.505 1.255 2.595 1.525 ;
        RECT  2.470 1.030 2.570 1.140 ;
        RECT  1.340 1.255 2.505 1.345 ;
        RECT  1.035 0.275 2.460 0.385 ;
        RECT  1.085 1.435 2.395 1.525 ;
        RECT  2.215 0.510 2.325 1.145 ;
        RECT  2.010 0.510 2.215 0.645 ;
        RECT  2.000 1.025 2.215 1.145 ;
        RECT  1.895 0.785 2.090 0.905 ;
        RECT  1.805 0.490 1.895 1.145 ;
        RECT  1.515 0.490 1.805 0.600 ;
        RECT  1.485 1.030 1.805 1.145 ;
        RECT  1.235 0.900 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFCNQD4

MACRO EDFD1
    CLASS CORE ;
    FOREIGN EDFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.220 0.300 5.350 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.455 4.950 1.285 ;
        RECT  4.705 0.455 4.850 0.625 ;
        RECT  4.705 1.115 4.850 1.285 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0661 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.710 1.750 0.910 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.165 5.400 0.165 ;
        RECT  3.070 0.490 3.220 0.595 ;
        RECT  2.980 -0.165 3.070 0.595 ;
        RECT  0.560 -0.165 2.980 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.155 1.635 5.400 1.965 ;
        RECT  2.985 1.435 3.155 1.965 ;
        RECT  0.475 1.635 2.985 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.040 0.275 5.130 1.505 ;
        RECT  3.985 0.275 5.040 0.365 ;
        RECT  3.390 1.410 5.040 1.505 ;
        RECT  4.615 0.750 4.750 0.920 ;
        RECT  4.525 0.455 4.615 1.320 ;
        RECT  4.225 0.455 4.525 0.575 ;
        RECT  4.390 1.215 4.525 1.320 ;
        RECT  4.345 0.750 4.435 1.125 ;
        RECT  4.005 1.035 4.345 1.125 ;
        RECT  4.115 0.455 4.225 0.920 ;
        RECT  3.915 0.600 4.005 1.320 ;
        RECT  3.895 0.275 3.985 0.490 ;
        RECT  3.805 0.600 3.915 0.690 ;
        RECT  3.525 1.230 3.915 1.320 ;
        RECT  3.715 0.295 3.805 0.690 ;
        RECT  3.690 0.830 3.800 1.135 ;
        RECT  3.575 0.295 3.715 0.415 ;
        RECT  3.620 0.830 3.690 0.940 ;
        RECT  3.510 0.525 3.620 0.940 ;
        RECT  3.420 0.275 3.445 0.445 ;
        RECT  3.325 0.275 3.420 1.165 ;
        RECT  3.300 1.255 3.390 1.505 ;
        RECT  2.845 0.995 3.325 1.165 ;
        RECT  1.340 1.255 3.300 1.345 ;
        RECT  2.690 0.710 3.235 0.880 ;
        RECT  2.600 0.305 2.690 1.145 ;
        RECT  2.490 1.035 2.600 1.145 ;
        RECT  1.035 0.275 2.490 0.385 ;
        RECT  1.085 1.435 2.410 1.525 ;
        RECT  2.230 0.510 2.340 1.145 ;
        RECT  2.025 0.510 2.230 0.645 ;
        RECT  2.030 1.025 2.230 1.145 ;
        RECT  1.930 0.785 2.105 0.905 ;
        RECT  1.840 0.490 1.930 1.145 ;
        RECT  1.530 0.490 1.840 0.600 ;
        RECT  1.500 1.030 1.840 1.145 ;
        RECT  1.230 0.915 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFD1

MACRO EDFD2
    CLASS CORE ;
    FOREIGN EDFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.350 0.455 5.525 0.595 ;
        RECT  5.350 1.180 5.525 1.320 ;
        RECT  5.250 0.455 5.350 1.320 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.455 5.150 1.320 ;
        RECT  4.835 0.455 5.050 0.595 ;
        RECT  4.815 1.110 5.050 1.320 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0661 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.710 1.750 0.910 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.060 -0.165 5.800 0.165 ;
        RECT  3.060 0.490 3.210 0.595 ;
        RECT  2.970 -0.165 3.060 0.595 ;
        RECT  0.560 -0.165 2.970 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.145 1.635 5.800 1.965 ;
        RECT  2.975 1.435 3.145 1.965 ;
        RECT  0.475 1.635 2.975 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.635 0.275 5.725 1.505 ;
        RECT  3.955 0.275 5.635 0.365 ;
        RECT  5.460 0.750 5.635 0.920 ;
        RECT  3.380 1.410 5.635 1.505 ;
        RECT  4.725 0.750 4.945 0.920 ;
        RECT  4.615 0.455 4.725 1.320 ;
        RECT  4.215 0.455 4.615 0.575 ;
        RECT  4.315 1.215 4.615 1.320 ;
        RECT  4.350 0.750 4.480 1.125 ;
        RECT  3.950 1.035 4.350 1.125 ;
        RECT  4.115 0.455 4.215 0.920 ;
        RECT  4.040 0.735 4.115 0.920 ;
        RECT  3.865 0.275 3.955 0.490 ;
        RECT  3.860 0.600 3.950 1.315 ;
        RECT  3.770 0.600 3.860 0.690 ;
        RECT  3.515 1.225 3.860 1.315 ;
        RECT  3.680 0.305 3.770 0.690 ;
        RECT  3.660 0.830 3.770 1.135 ;
        RECT  3.565 0.305 3.680 0.415 ;
        RECT  3.590 0.830 3.660 0.940 ;
        RECT  3.500 0.525 3.590 0.940 ;
        RECT  3.410 0.275 3.475 0.385 ;
        RECT  3.315 0.275 3.410 1.165 ;
        RECT  3.290 1.255 3.380 1.505 ;
        RECT  3.285 0.275 3.315 0.385 ;
        RECT  2.835 0.995 3.315 1.165 ;
        RECT  1.340 1.255 3.290 1.345 ;
        RECT  2.680 0.710 3.225 0.880 ;
        RECT  2.590 0.305 2.680 1.145 ;
        RECT  2.480 1.035 2.590 1.145 ;
        RECT  1.035 0.275 2.480 0.385 ;
        RECT  1.085 1.435 2.400 1.525 ;
        RECT  2.220 0.510 2.330 1.145 ;
        RECT  2.025 0.510 2.220 0.645 ;
        RECT  2.020 1.025 2.220 1.145 ;
        RECT  1.930 0.785 2.105 0.905 ;
        RECT  1.840 0.490 1.930 1.145 ;
        RECT  1.530 0.490 1.840 0.600 ;
        RECT  1.500 1.030 1.840 1.145 ;
        RECT  1.230 0.915 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFD2

MACRO EDFD4
    CLASS CORE ;
    FOREIGN EDFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.295 7.080 0.665 ;
        RECT  6.850 1.080 7.080 1.450 ;
        RECT  6.550 0.295 6.850 1.450 ;
        RECT  6.415 0.295 6.550 0.665 ;
        RECT  6.410 1.080 6.550 1.450 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.455 6.100 0.635 ;
        RECT  6.050 1.075 6.100 1.300 ;
        RECT  5.750 0.455 6.050 1.300 ;
        RECT  5.385 0.455 5.750 0.635 ;
        RECT  5.385 1.055 5.750 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0643 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.710 1.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.320 -0.165 7.400 0.165 ;
        RECT  7.190 -0.165 7.320 0.685 ;
        RECT  3.120 -0.165 7.190 0.165 ;
        RECT  3.120 0.490 3.215 0.595 ;
        RECT  3.030 -0.165 3.120 0.595 ;
        RECT  0.560 -0.165 3.030 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.315 1.635 7.400 1.965 ;
        RECT  7.195 1.015 7.315 1.965 ;
        RECT  3.205 1.635 7.195 1.965 ;
        RECT  3.035 1.435 3.205 1.965 ;
        RECT  0.475 1.635 3.035 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.950 0.295 7.080 0.665 ;
        RECT  6.950 1.080 7.080 1.450 ;
        RECT  6.415 0.295 6.450 0.665 ;
        RECT  6.410 1.080 6.450 1.450 ;
        RECT  5.385 0.455 5.650 0.635 ;
        RECT  5.385 1.055 5.650 1.300 ;
        RECT  6.300 0.770 6.440 0.940 ;
        RECT  6.210 0.275 6.300 1.505 ;
        RECT  4.525 0.275 6.210 0.365 ;
        RECT  4.525 1.410 6.210 1.505 ;
        RECT  5.275 0.765 5.620 0.910 ;
        RECT  5.165 0.455 5.275 1.320 ;
        RECT  4.765 0.455 5.165 0.575 ;
        RECT  4.865 1.215 5.165 1.320 ;
        RECT  4.900 0.750 5.030 1.125 ;
        RECT  4.150 1.035 4.900 1.125 ;
        RECT  4.665 0.455 4.765 0.900 ;
        RECT  4.345 0.775 4.665 0.900 ;
        RECT  4.395 0.275 4.525 0.645 ;
        RECT  4.395 1.245 4.525 1.505 ;
        RECT  3.990 0.275 4.395 0.365 ;
        RECT  3.440 1.410 4.395 1.505 ;
        RECT  4.030 0.600 4.150 1.320 ;
        RECT  3.790 0.600 4.030 0.690 ;
        RECT  3.575 1.230 4.030 1.320 ;
        RECT  3.880 0.275 3.990 0.470 ;
        RECT  3.740 0.830 3.860 1.140 ;
        RECT  3.700 0.310 3.790 0.690 ;
        RECT  3.610 0.830 3.740 0.940 ;
        RECT  3.590 0.310 3.700 0.420 ;
        RECT  3.520 0.530 3.610 0.940 ;
        RECT  3.430 0.275 3.500 0.385 ;
        RECT  3.430 1.035 3.490 1.165 ;
        RECT  3.350 1.255 3.440 1.505 ;
        RECT  3.340 0.275 3.430 1.165 ;
        RECT  1.340 1.255 3.350 1.345 ;
        RECT  3.330 0.275 3.340 0.595 ;
        RECT  2.895 0.995 3.340 1.165 ;
        RECT  2.740 0.710 3.250 0.880 ;
        RECT  2.595 0.305 2.740 1.145 ;
        RECT  2.540 1.035 2.595 1.145 ;
        RECT  1.035 0.275 2.485 0.385 ;
        RECT  1.085 1.435 2.445 1.525 ;
        RECT  2.260 0.510 2.360 1.145 ;
        RECT  2.045 0.510 2.260 0.645 ;
        RECT  2.035 1.025 2.260 1.145 ;
        RECT  1.945 0.750 2.030 0.920 ;
        RECT  1.855 0.490 1.945 1.145 ;
        RECT  1.550 0.490 1.855 0.600 ;
        RECT  1.520 1.030 1.855 1.145 ;
        RECT  1.235 0.900 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFD4

MACRO EDFKCND1
    CLASS CORE ;
    FOREIGN EDFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.285 5.750 1.515 ;
        RECT  5.625 0.285 5.650 0.665 ;
        RECT  5.625 1.015 5.650 1.515 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.260 0.455 5.350 1.300 ;
        RECT  5.075 0.455 5.260 0.690 ;
        RECT  5.075 1.055 5.260 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.120 ;
        RECT  0.180 0.800 0.245 1.005 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.935 0.965 1.045 ;
        RECT  0.650 0.935 0.755 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.475 -0.165 5.800 0.165 ;
        RECT  3.475 0.490 3.570 0.595 ;
        RECT  3.385 -0.165 3.475 0.595 ;
        RECT  0.555 -0.165 3.385 0.165 ;
        RECT  0.465 -0.165 0.555 0.395 ;
        RECT  0.000 -0.165 0.465 0.165 ;
        RECT  0.285 0.285 0.465 0.395 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.635 5.800 1.965 ;
        RECT  3.390 1.435 3.560 1.965 ;
        RECT  0.495 1.635 3.390 1.965 ;
        RECT  0.305 1.395 0.495 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.535 0.770 5.550 0.940 ;
        RECT  5.445 0.275 5.535 1.505 ;
        RECT  4.370 0.275 5.445 0.365 ;
        RECT  3.795 1.410 5.445 1.505 ;
        RECT  4.985 0.780 5.095 0.900 ;
        RECT  4.875 0.455 4.985 1.320 ;
        RECT  4.555 0.455 4.875 0.575 ;
        RECT  4.740 1.215 4.875 1.320 ;
        RECT  4.675 0.750 4.785 1.125 ;
        RECT  4.375 1.035 4.675 1.125 ;
        RECT  4.465 0.455 4.555 0.920 ;
        RECT  4.285 0.600 4.375 1.320 ;
        RECT  4.260 0.275 4.370 0.460 ;
        RECT  4.145 0.600 4.285 0.690 ;
        RECT  3.930 1.230 4.285 1.320 ;
        RECT  4.075 0.830 4.195 1.140 ;
        RECT  4.055 0.310 4.145 0.690 ;
        RECT  3.965 0.830 4.075 0.940 ;
        RECT  3.945 0.310 4.055 0.420 ;
        RECT  3.875 0.530 3.965 0.940 ;
        RECT  3.785 0.275 3.855 0.385 ;
        RECT  3.785 1.035 3.845 1.140 ;
        RECT  3.705 1.230 3.795 1.505 ;
        RECT  3.695 0.275 3.785 1.140 ;
        RECT  1.475 1.230 3.705 1.320 ;
        RECT  3.685 0.275 3.695 0.595 ;
        RECT  3.250 0.995 3.695 1.140 ;
        RECT  3.095 0.725 3.605 0.895 ;
        RECT  2.950 0.305 3.095 1.140 ;
        RECT  2.875 1.015 2.950 1.140 ;
        RECT  1.150 0.275 2.840 0.385 ;
        RECT  1.075 1.410 2.800 1.505 ;
        RECT  2.615 0.525 2.715 1.140 ;
        RECT  2.420 0.525 2.615 0.640 ;
        RECT  2.420 1.025 2.615 1.140 ;
        RECT  2.330 0.750 2.385 0.920 ;
        RECT  2.240 0.510 2.330 1.140 ;
        RECT  1.900 0.510 2.240 0.620 ;
        RECT  1.900 1.030 2.240 1.140 ;
        RECT  1.385 0.800 1.475 1.320 ;
        RECT  1.095 0.755 1.225 0.965 ;
        RECT  0.980 0.275 1.150 0.655 ;
        RECT  0.540 0.755 1.095 0.845 ;
        RECT  0.945 1.250 1.075 1.505 ;
        RECT  0.450 0.490 0.540 1.305 ;
        RECT  0.185 0.490 0.450 0.580 ;
        RECT  0.185 1.215 0.450 1.305 ;
        RECT  0.075 0.295 0.185 0.580 ;
        RECT  0.075 1.215 0.185 1.505 ;
    END
END EDFKCND1

MACRO EDFKCND2
    CLASS CORE ;
    FOREIGN EDFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.830 0.285 5.950 1.515 ;
        RECT  5.775 0.285 5.830 0.690 ;
        RECT  5.775 1.015 5.830 1.515 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.370 0.455 5.460 1.300 ;
        RECT  5.235 0.455 5.370 0.690 ;
        RECT  5.235 1.055 5.370 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.120 ;
        RECT  0.180 0.800 0.245 1.005 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.935 0.965 1.045 ;
        RECT  0.650 0.935 0.755 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.475 -0.165 6.200 0.165 ;
        RECT  3.475 0.490 3.570 0.595 ;
        RECT  3.385 -0.165 3.475 0.595 ;
        RECT  0.555 -0.165 3.385 0.165 ;
        RECT  0.465 -0.165 0.555 0.395 ;
        RECT  0.000 -0.165 0.465 0.165 ;
        RECT  0.285 0.285 0.465 0.395 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.635 6.200 1.965 ;
        RECT  3.390 1.435 3.560 1.965 ;
        RECT  0.495 1.635 3.390 1.965 ;
        RECT  0.305 1.395 0.495 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.665 0.770 5.700 0.940 ;
        RECT  5.550 0.275 5.665 1.505 ;
        RECT  4.345 0.275 5.550 0.365 ;
        RECT  3.795 1.410 5.550 1.505 ;
        RECT  5.125 0.780 5.280 0.900 ;
        RECT  5.015 0.455 5.125 1.320 ;
        RECT  4.530 0.455 5.015 0.575 ;
        RECT  4.715 1.215 5.015 1.320 ;
        RECT  4.750 0.750 4.880 1.125 ;
        RECT  4.350 1.035 4.750 1.125 ;
        RECT  4.440 0.455 4.530 0.920 ;
        RECT  4.260 0.600 4.350 1.320 ;
        RECT  4.235 0.275 4.345 0.460 ;
        RECT  4.145 0.600 4.260 0.690 ;
        RECT  3.930 1.230 4.260 1.320 ;
        RECT  4.060 0.830 4.170 1.140 ;
        RECT  4.055 0.310 4.145 0.690 ;
        RECT  3.965 0.830 4.060 0.940 ;
        RECT  3.945 0.310 4.055 0.420 ;
        RECT  3.875 0.530 3.965 0.940 ;
        RECT  3.785 0.275 3.855 0.385 ;
        RECT  3.785 1.035 3.845 1.140 ;
        RECT  3.705 1.230 3.795 1.505 ;
        RECT  3.695 0.275 3.785 1.140 ;
        RECT  1.475 1.230 3.705 1.320 ;
        RECT  3.685 0.275 3.695 0.595 ;
        RECT  3.250 0.995 3.695 1.140 ;
        RECT  3.095 0.725 3.605 0.895 ;
        RECT  2.950 0.305 3.095 1.140 ;
        RECT  2.875 1.015 2.950 1.140 ;
        RECT  1.150 0.275 2.840 0.385 ;
        RECT  1.075 1.410 2.800 1.505 ;
        RECT  2.615 0.525 2.715 1.140 ;
        RECT  2.420 0.525 2.615 0.640 ;
        RECT  2.420 1.025 2.615 1.140 ;
        RECT  2.330 0.750 2.385 0.920 ;
        RECT  2.240 0.510 2.330 1.140 ;
        RECT  1.900 0.510 2.240 0.620 ;
        RECT  1.900 1.030 2.240 1.140 ;
        RECT  1.385 0.800 1.475 1.320 ;
        RECT  1.095 0.755 1.225 0.965 ;
        RECT  0.980 0.275 1.150 0.655 ;
        RECT  0.540 0.755 1.095 0.845 ;
        RECT  0.945 1.250 1.075 1.505 ;
        RECT  0.450 0.490 0.540 1.305 ;
        RECT  0.185 0.490 0.450 0.580 ;
        RECT  0.185 1.215 0.450 1.305 ;
        RECT  0.075 0.295 0.185 0.580 ;
        RECT  0.075 1.215 0.185 1.505 ;
    END
END EDFKCND2

MACRO EDFKCND4
    CLASS CORE ;
    FOREIGN EDFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.295 7.480 0.665 ;
        RECT  7.250 1.080 7.480 1.450 ;
        RECT  6.950 0.295 7.250 1.450 ;
        RECT  6.815 0.295 6.950 0.665 ;
        RECT  6.810 1.080 6.950 1.450 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.455 6.500 0.635 ;
        RECT  6.450 1.075 6.500 1.300 ;
        RECT  6.150 0.455 6.450 1.300 ;
        RECT  5.785 0.455 6.150 0.635 ;
        RECT  5.785 1.055 6.150 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.120 ;
        RECT  0.180 0.800 0.245 1.005 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.935 0.965 1.045 ;
        RECT  0.650 0.935 0.755 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.160 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.720 -0.165 7.800 0.165 ;
        RECT  7.590 -0.165 7.720 0.685 ;
        RECT  3.520 -0.165 7.590 0.165 ;
        RECT  3.520 0.490 3.615 0.595 ;
        RECT  3.430 -0.165 3.520 0.595 ;
        RECT  0.555 -0.165 3.430 0.165 ;
        RECT  0.465 -0.165 0.555 0.395 ;
        RECT  0.000 -0.165 0.465 0.165 ;
        RECT  0.285 0.285 0.465 0.395 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.715 1.635 7.800 1.965 ;
        RECT  7.595 1.015 7.715 1.965 ;
        RECT  3.605 1.635 7.595 1.965 ;
        RECT  3.435 1.435 3.605 1.965 ;
        RECT  0.495 1.635 3.435 1.965 ;
        RECT  0.305 1.395 0.495 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.350 0.295 7.480 0.665 ;
        RECT  7.350 1.080 7.480 1.450 ;
        RECT  6.815 0.295 6.850 0.665 ;
        RECT  6.810 1.080 6.850 1.450 ;
        RECT  5.785 0.455 6.050 0.635 ;
        RECT  5.785 1.055 6.050 1.300 ;
        RECT  6.700 0.770 6.840 0.940 ;
        RECT  6.610 0.275 6.700 1.505 ;
        RECT  4.925 0.275 6.610 0.365 ;
        RECT  4.925 1.410 6.610 1.505 ;
        RECT  5.675 0.765 6.020 0.910 ;
        RECT  5.565 0.455 5.675 1.320 ;
        RECT  5.165 0.455 5.565 0.575 ;
        RECT  5.265 1.215 5.565 1.320 ;
        RECT  5.300 0.750 5.430 1.125 ;
        RECT  4.530 1.035 5.300 1.125 ;
        RECT  5.065 0.455 5.165 0.900 ;
        RECT  4.745 0.775 5.065 0.900 ;
        RECT  4.795 0.275 4.925 0.645 ;
        RECT  4.795 1.245 4.925 1.505 ;
        RECT  4.390 0.275 4.795 0.365 ;
        RECT  3.840 1.410 4.795 1.505 ;
        RECT  4.430 0.600 4.530 1.320 ;
        RECT  4.190 0.600 4.430 0.690 ;
        RECT  3.975 1.230 4.430 1.320 ;
        RECT  4.280 0.275 4.390 0.460 ;
        RECT  4.150 0.830 4.270 1.140 ;
        RECT  4.100 0.305 4.190 0.690 ;
        RECT  4.010 0.830 4.150 0.940 ;
        RECT  3.990 0.305 4.100 0.415 ;
        RECT  3.920 0.530 4.010 0.940 ;
        RECT  3.830 0.275 3.900 0.385 ;
        RECT  3.830 1.035 3.890 1.140 ;
        RECT  3.750 1.230 3.840 1.505 ;
        RECT  3.740 0.275 3.830 1.140 ;
        RECT  1.475 1.230 3.750 1.320 ;
        RECT  3.730 0.275 3.740 0.595 ;
        RECT  3.295 0.995 3.740 1.140 ;
        RECT  3.140 0.725 3.650 0.895 ;
        RECT  2.995 0.305 3.140 1.140 ;
        RECT  2.920 1.015 2.995 1.140 ;
        RECT  1.150 0.275 2.885 0.385 ;
        RECT  1.075 1.410 2.845 1.505 ;
        RECT  2.660 0.510 2.760 1.140 ;
        RECT  2.445 0.510 2.660 0.645 ;
        RECT  2.435 1.025 2.660 1.140 ;
        RECT  2.345 0.750 2.430 0.920 ;
        RECT  2.255 0.490 2.345 1.140 ;
        RECT  1.965 0.490 2.255 0.600 ;
        RECT  1.890 1.030 2.255 1.140 ;
        RECT  1.385 0.800 1.475 1.320 ;
        RECT  1.095 0.755 1.225 0.955 ;
        RECT  0.980 0.275 1.150 0.655 ;
        RECT  0.540 0.755 1.095 0.845 ;
        RECT  0.945 1.250 1.075 1.505 ;
        RECT  0.450 0.490 0.540 1.305 ;
        RECT  0.185 0.490 0.450 0.580 ;
        RECT  0.185 1.215 0.450 1.305 ;
        RECT  0.075 0.295 0.185 0.580 ;
        RECT  0.075 1.215 0.185 1.505 ;
    END
END EDFKCND4

MACRO EDFKCNQD1
    CLASS CORE ;
    FOREIGN EDFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.510 5.350 1.290 ;
        RECT  5.085 0.510 5.250 0.690 ;
        RECT  5.085 1.110 5.250 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0775 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.120 ;
        RECT  0.180 0.800 0.245 1.005 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.935 0.965 1.045 ;
        RECT  0.650 0.935 0.750 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.505 -0.165 5.600 0.165 ;
        RECT  3.505 0.490 3.600 0.595 ;
        RECT  3.415 -0.165 3.505 0.595 ;
        RECT  0.555 -0.165 3.415 0.165 ;
        RECT  0.465 -0.165 0.555 0.395 ;
        RECT  0.000 -0.165 0.465 0.165 ;
        RECT  0.285 0.285 0.465 0.395 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.635 5.600 1.965 ;
        RECT  3.420 1.435 3.590 1.965 ;
        RECT  0.495 1.635 3.420 1.965 ;
        RECT  0.310 1.395 0.495 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.440 0.275 5.550 1.505 ;
        RECT  4.380 0.275 5.440 0.365 ;
        RECT  3.825 1.410 5.440 1.505 ;
        RECT  4.995 0.780 5.145 0.910 ;
        RECT  4.905 0.455 4.995 1.320 ;
        RECT  4.605 0.455 4.905 0.565 ;
        RECT  4.770 1.210 4.905 1.320 ;
        RECT  4.725 0.725 4.815 1.115 ;
        RECT  4.405 1.015 4.725 1.115 ;
        RECT  4.495 0.455 4.605 0.920 ;
        RECT  4.315 0.600 4.405 1.320 ;
        RECT  4.270 0.275 4.380 0.460 ;
        RECT  4.175 0.600 4.315 0.690 ;
        RECT  3.960 1.230 4.315 1.320 ;
        RECT  4.115 0.830 4.225 1.140 ;
        RECT  4.085 0.310 4.175 0.690 ;
        RECT  3.995 0.830 4.115 0.940 ;
        RECT  3.975 0.310 4.085 0.420 ;
        RECT  3.905 0.530 3.995 0.940 ;
        RECT  3.815 0.275 3.885 0.385 ;
        RECT  3.815 1.035 3.875 1.125 ;
        RECT  3.735 1.215 3.825 1.505 ;
        RECT  3.725 0.275 3.815 1.125 ;
        RECT  1.495 1.215 3.735 1.305 ;
        RECT  3.715 0.275 3.725 0.595 ;
        RECT  3.280 0.995 3.725 1.125 ;
        RECT  3.125 0.725 3.635 0.895 ;
        RECT  2.980 0.305 3.125 1.125 ;
        RECT  2.905 1.000 2.980 1.125 ;
        RECT  1.150 0.275 2.870 0.385 ;
        RECT  1.070 1.395 2.820 1.525 ;
        RECT  2.635 0.475 2.735 1.125 ;
        RECT  2.445 0.475 2.635 0.645 ;
        RECT  2.445 1.010 2.635 1.125 ;
        RECT  2.355 0.750 2.385 0.920 ;
        RECT  2.265 0.510 2.355 1.125 ;
        RECT  1.875 0.510 2.265 0.620 ;
        RECT  1.865 1.015 2.265 1.125 ;
        RECT  1.385 0.780 1.495 1.305 ;
        RECT  1.095 0.755 1.225 0.965 ;
        RECT  0.980 0.275 1.150 0.655 ;
        RECT  0.540 0.755 1.095 0.845 ;
        RECT  0.955 1.250 1.070 1.525 ;
        RECT  0.450 0.490 0.540 1.305 ;
        RECT  0.185 0.490 0.450 0.580 ;
        RECT  0.185 1.215 0.450 1.305 ;
        RECT  0.075 0.295 0.185 0.580 ;
        RECT  0.075 1.215 0.185 1.505 ;
    END
END EDFKCNQD1

MACRO EDFKCNQD2
    CLASS CORE ;
    FOREIGN EDFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.455 5.550 1.300 ;
        RECT  5.255 0.455 5.450 0.635 ;
        RECT  5.250 1.055 5.450 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.120 ;
        RECT  0.180 0.800 0.245 1.005 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.935 0.965 1.045 ;
        RECT  0.650 0.935 0.750 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.730 2.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0527 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.470 -0.165 5.800 0.165 ;
        RECT  3.470 0.490 3.565 0.595 ;
        RECT  3.380 -0.165 3.470 0.595 ;
        RECT  0.555 -0.165 3.380 0.165 ;
        RECT  0.465 -0.165 0.555 0.395 ;
        RECT  0.000 -0.165 0.465 0.165 ;
        RECT  0.285 0.285 0.465 0.395 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.555 1.635 5.800 1.965 ;
        RECT  3.385 1.435 3.555 1.965 ;
        RECT  0.495 1.635 3.385 1.965 ;
        RECT  0.310 1.395 0.495 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.650 0.275 5.750 1.505 ;
        RECT  4.365 0.275 5.650 0.365 ;
        RECT  3.790 1.410 5.650 1.505 ;
        RECT  5.145 0.765 5.360 0.910 ;
        RECT  5.035 0.455 5.145 1.320 ;
        RECT  4.625 0.455 5.035 0.575 ;
        RECT  4.735 1.215 5.035 1.320 ;
        RECT  4.770 0.750 4.900 1.125 ;
        RECT  4.370 1.035 4.770 1.125 ;
        RECT  4.525 0.455 4.625 0.920 ;
        RECT  4.460 0.750 4.525 0.920 ;
        RECT  4.280 0.600 4.370 1.320 ;
        RECT  4.255 0.275 4.365 0.460 ;
        RECT  4.140 0.600 4.280 0.690 ;
        RECT  3.925 1.230 4.280 1.320 ;
        RECT  4.080 0.830 4.190 1.140 ;
        RECT  4.050 0.310 4.140 0.690 ;
        RECT  3.960 0.830 4.080 0.940 ;
        RECT  3.940 0.310 4.050 0.420 ;
        RECT  3.870 0.530 3.960 0.940 ;
        RECT  3.780 0.275 3.850 0.385 ;
        RECT  3.780 1.035 3.840 1.140 ;
        RECT  3.700 1.230 3.790 1.505 ;
        RECT  3.690 0.275 3.780 1.140 ;
        RECT  1.485 1.230 3.700 1.320 ;
        RECT  3.680 0.275 3.690 0.595 ;
        RECT  3.245 0.995 3.690 1.140 ;
        RECT  3.090 0.710 3.600 0.880 ;
        RECT  2.945 0.305 3.090 1.140 ;
        RECT  2.870 1.015 2.945 1.140 ;
        RECT  1.150 0.275 2.835 0.385 ;
        RECT  1.895 1.410 2.795 1.505 ;
        RECT  2.610 0.475 2.710 1.140 ;
        RECT  2.435 0.475 2.610 0.645 ;
        RECT  2.420 1.025 2.610 1.140 ;
        RECT  2.330 0.750 2.380 0.920 ;
        RECT  2.240 0.490 2.330 1.140 ;
        RECT  1.915 0.490 2.240 0.600 ;
        RECT  1.840 1.030 2.240 1.140 ;
        RECT  1.725 1.410 1.895 1.515 ;
        RECT  1.070 1.410 1.725 1.505 ;
        RECT  1.370 0.780 1.485 1.320 ;
        RECT  1.095 0.755 1.225 0.955 ;
        RECT  0.980 0.275 1.150 0.655 ;
        RECT  0.540 0.755 1.095 0.845 ;
        RECT  0.955 1.250 1.070 1.505 ;
        RECT  0.450 0.490 0.540 1.305 ;
        RECT  0.185 0.490 0.450 0.580 ;
        RECT  0.185 1.215 0.450 1.305 ;
        RECT  0.075 0.295 0.185 0.580 ;
        RECT  0.075 1.215 0.185 1.505 ;
    END
END EDFKCNQD2

MACRO EDFKCNQD4
    CLASS CORE ;
    FOREIGN EDFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.455 5.905 0.635 ;
        RECT  5.850 1.075 5.905 1.300 ;
        RECT  5.550 0.455 5.850 1.300 ;
        RECT  5.230 0.455 5.550 0.635 ;
        RECT  5.230 1.055 5.550 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.120 ;
        RECT  0.180 0.800 0.245 1.005 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.935 0.965 1.045 ;
        RECT  0.650 0.935 0.755 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.730 2.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.750 1.110 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.470 -0.165 6.200 0.165 ;
        RECT  3.470 0.490 3.565 0.595 ;
        RECT  3.380 -0.165 3.470 0.595 ;
        RECT  0.555 -0.165 3.380 0.165 ;
        RECT  0.465 -0.165 0.555 0.395 ;
        RECT  0.000 -0.165 0.465 0.165 ;
        RECT  0.285 0.285 0.465 0.395 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.555 1.635 6.200 1.965 ;
        RECT  3.385 1.435 3.555 1.965 ;
        RECT  0.495 1.635 3.385 1.965 ;
        RECT  0.305 1.395 0.495 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.230 0.455 5.450 0.635 ;
        RECT  5.230 1.055 5.450 1.300 ;
        RECT  6.015 0.275 6.115 1.505 ;
        RECT  4.340 0.275 6.015 0.365 ;
        RECT  3.790 1.410 6.015 1.505 ;
        RECT  5.120 0.765 5.445 0.910 ;
        RECT  5.010 0.455 5.120 1.320 ;
        RECT  4.600 0.455 5.010 0.575 ;
        RECT  4.710 1.215 5.010 1.320 ;
        RECT  4.745 0.750 4.875 1.125 ;
        RECT  4.345 1.035 4.745 1.125 ;
        RECT  4.500 0.455 4.600 0.920 ;
        RECT  4.435 0.750 4.500 0.920 ;
        RECT  4.255 0.600 4.345 1.320 ;
        RECT  4.230 0.275 4.340 0.460 ;
        RECT  4.140 0.600 4.255 0.690 ;
        RECT  3.925 1.230 4.255 1.320 ;
        RECT  4.055 0.830 4.165 1.140 ;
        RECT  4.050 0.310 4.140 0.690 ;
        RECT  3.960 0.830 4.055 0.940 ;
        RECT  3.940 0.310 4.050 0.420 ;
        RECT  3.870 0.530 3.960 0.940 ;
        RECT  3.780 0.275 3.850 0.385 ;
        RECT  3.780 1.035 3.840 1.140 ;
        RECT  3.700 1.230 3.790 1.505 ;
        RECT  3.690 0.275 3.780 1.140 ;
        RECT  1.485 1.230 3.700 1.320 ;
        RECT  3.680 0.275 3.690 0.595 ;
        RECT  3.245 0.995 3.690 1.140 ;
        RECT  3.090 0.725 3.600 0.895 ;
        RECT  2.945 0.305 3.090 1.140 ;
        RECT  2.870 1.015 2.945 1.140 ;
        RECT  1.150 0.275 2.835 0.385 ;
        RECT  1.075 1.410 2.795 1.505 ;
        RECT  2.610 0.475 2.710 1.140 ;
        RECT  2.435 0.475 2.610 0.645 ;
        RECT  2.420 1.025 2.610 1.140 ;
        RECT  2.330 0.750 2.380 0.920 ;
        RECT  2.240 0.490 2.330 1.140 ;
        RECT  1.915 0.490 2.240 0.600 ;
        RECT  1.840 1.030 2.240 1.140 ;
        RECT  1.365 0.780 1.485 1.320 ;
        RECT  1.095 0.755 1.225 0.955 ;
        RECT  0.980 0.275 1.150 0.655 ;
        RECT  0.540 0.755 1.095 0.845 ;
        RECT  0.945 1.250 1.075 1.505 ;
        RECT  0.450 0.490 0.540 1.305 ;
        RECT  0.185 0.490 0.450 0.580 ;
        RECT  0.185 1.215 0.450 1.305 ;
        RECT  0.075 0.295 0.185 0.580 ;
        RECT  0.075 1.215 0.185 1.505 ;
    END
END EDFKCNQD4

MACRO EDFQD1
    CLASS CORE ;
    FOREIGN EDFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.455 4.950 1.320 ;
        RECT  4.650 0.455 4.850 0.595 ;
        RECT  4.650 1.110 4.850 1.320 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0643 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.800 1.710 0.910 ;
        RECT  1.435 0.690 1.550 0.910 ;
        RECT  1.370 0.690 1.435 0.790 ;
        RECT  1.245 0.510 1.370 0.790 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.060 -0.165 5.200 0.165 ;
        RECT  3.060 0.490 3.210 0.595 ;
        RECT  2.970 -0.165 3.060 0.595 ;
        RECT  0.560 -0.165 2.970 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.145 1.635 5.200 1.965 ;
        RECT  2.975 1.435 3.145 1.965 ;
        RECT  0.475 1.635 2.975 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.040 0.275 5.130 1.505 ;
        RECT  3.955 0.275 5.040 0.365 ;
        RECT  3.380 1.410 5.040 1.505 ;
        RECT  4.560 0.750 4.750 0.920 ;
        RECT  4.460 0.455 4.560 1.320 ;
        RECT  4.160 0.455 4.460 0.575 ;
        RECT  4.355 1.215 4.460 1.320 ;
        RECT  4.250 0.750 4.370 1.125 ;
        RECT  3.960 1.035 4.250 1.125 ;
        RECT  4.050 0.455 4.160 0.920 ;
        RECT  3.870 0.600 3.960 1.320 ;
        RECT  3.865 0.275 3.955 0.490 ;
        RECT  3.770 0.600 3.870 0.690 ;
        RECT  3.515 1.230 3.870 1.320 ;
        RECT  3.670 0.830 3.780 1.140 ;
        RECT  3.680 0.310 3.770 0.690 ;
        RECT  3.565 0.310 3.680 0.420 ;
        RECT  3.590 0.830 3.670 0.940 ;
        RECT  3.500 0.530 3.590 0.940 ;
        RECT  3.410 0.275 3.475 0.385 ;
        RECT  3.315 0.275 3.410 1.165 ;
        RECT  3.290 1.255 3.380 1.505 ;
        RECT  3.285 0.275 3.315 0.385 ;
        RECT  2.835 0.995 3.315 1.165 ;
        RECT  1.340 1.255 3.290 1.345 ;
        RECT  2.680 0.725 3.225 0.895 ;
        RECT  2.590 0.305 2.680 1.145 ;
        RECT  2.480 1.035 2.590 1.145 ;
        RECT  1.035 0.275 2.480 0.385 ;
        RECT  1.085 1.435 2.385 1.525 ;
        RECT  2.225 0.510 2.335 1.145 ;
        RECT  2.035 0.510 2.225 0.645 ;
        RECT  2.015 1.025 2.225 1.145 ;
        RECT  1.910 0.785 2.105 0.905 ;
        RECT  1.820 0.490 1.910 1.145 ;
        RECT  1.540 0.490 1.820 0.600 ;
        RECT  1.500 1.030 1.820 1.145 ;
        RECT  1.235 0.900 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFQD1

MACRO EDFQD2
    CLASS CORE ;
    FOREIGN EDFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1780 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.455 5.150 1.320 ;
        RECT  4.895 0.455 5.050 0.595 ;
        RECT  4.875 1.180 5.050 1.320 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0643 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.800 1.710 0.910 ;
        RECT  1.435 0.690 1.550 0.910 ;
        RECT  1.370 0.690 1.435 0.790 ;
        RECT  1.245 0.510 1.370 0.790 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.060 -0.165 5.400 0.165 ;
        RECT  3.060 0.490 3.210 0.595 ;
        RECT  2.970 -0.165 3.060 0.595 ;
        RECT  0.560 -0.165 2.970 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.145 1.635 5.400 1.965 ;
        RECT  2.975 1.435 3.145 1.965 ;
        RECT  0.475 1.635 2.975 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.240 0.275 5.340 1.505 ;
        RECT  3.980 0.275 5.240 0.365 ;
        RECT  3.380 1.410 5.240 1.505 ;
        RECT  4.785 0.750 4.830 0.920 ;
        RECT  4.675 0.455 4.785 1.320 ;
        RECT  4.230 0.455 4.675 0.575 ;
        RECT  4.345 1.215 4.675 1.320 ;
        RECT  4.380 0.750 4.510 1.125 ;
        RECT  3.960 1.035 4.380 1.125 ;
        RECT  4.140 0.455 4.230 0.920 ;
        RECT  4.050 0.735 4.140 0.920 ;
        RECT  3.890 0.275 3.980 0.490 ;
        RECT  3.870 0.600 3.960 1.320 ;
        RECT  3.770 0.600 3.870 0.690 ;
        RECT  3.515 1.230 3.870 1.320 ;
        RECT  3.670 0.830 3.780 1.140 ;
        RECT  3.680 0.310 3.770 0.690 ;
        RECT  3.565 0.310 3.680 0.420 ;
        RECT  3.590 0.830 3.670 0.940 ;
        RECT  3.500 0.530 3.590 0.940 ;
        RECT  3.410 0.275 3.475 0.420 ;
        RECT  3.315 0.275 3.410 1.165 ;
        RECT  3.290 1.255 3.380 1.505 ;
        RECT  3.285 0.275 3.315 0.385 ;
        RECT  2.835 0.995 3.315 1.165 ;
        RECT  1.340 1.255 3.290 1.345 ;
        RECT  2.680 0.725 3.225 0.895 ;
        RECT  2.590 0.305 2.680 1.145 ;
        RECT  2.480 1.035 2.590 1.145 ;
        RECT  1.035 0.275 2.480 0.385 ;
        RECT  1.085 1.435 2.385 1.525 ;
        RECT  2.225 0.510 2.335 1.145 ;
        RECT  2.035 0.510 2.225 0.645 ;
        RECT  2.015 1.025 2.225 1.145 ;
        RECT  1.910 0.785 2.105 0.905 ;
        RECT  1.820 0.490 1.910 1.145 ;
        RECT  1.540 0.490 1.820 0.600 ;
        RECT  1.500 1.030 1.820 1.145 ;
        RECT  1.235 0.900 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFQD2

MACRO EDFQD4
    CLASS CORE ;
    FOREIGN EDFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.475 5.660 0.690 ;
        RECT  5.450 1.055 5.660 1.300 ;
        RECT  5.150 0.475 5.450 1.300 ;
        RECT  4.945 0.475 5.150 0.665 ;
        RECT  4.945 1.055 5.150 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0643 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.750 0.590 0.920 ;
        RECT  0.450 0.510 0.560 0.920 ;
        RECT  0.400 0.510 0.450 0.600 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.710 1.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.120 -0.165 6.000 0.165 ;
        RECT  3.120 0.490 3.215 0.595 ;
        RECT  3.030 -0.165 3.120 0.595 ;
        RECT  0.560 -0.165 3.030 0.165 ;
        RECT  0.440 -0.165 0.560 0.410 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        RECT  0.305 0.300 0.440 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.205 1.635 6.000 1.965 ;
        RECT  3.035 1.435 3.205 1.965 ;
        RECT  0.475 1.635 3.035 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.550 0.475 5.660 0.690 ;
        RECT  5.550 1.055 5.660 1.300 ;
        RECT  4.945 0.475 5.050 0.665 ;
        RECT  4.945 1.055 5.050 1.300 ;
        RECT  5.770 0.275 5.870 1.505 ;
        RECT  3.990 0.275 5.770 0.365 ;
        RECT  3.440 1.410 5.770 1.505 ;
        RECT  4.835 0.765 5.040 0.910 ;
        RECT  4.700 0.455 4.835 1.320 ;
        RECT  4.245 0.455 4.700 0.575 ;
        RECT  4.400 1.215 4.700 1.320 ;
        RECT  4.435 0.750 4.565 1.125 ;
        RECT  4.020 1.035 4.435 1.125 ;
        RECT  4.125 0.455 4.245 0.920 ;
        RECT  3.930 0.600 4.020 1.320 ;
        RECT  3.880 0.275 3.990 0.470 ;
        RECT  3.790 0.600 3.930 0.690 ;
        RECT  3.575 1.230 3.930 1.320 ;
        RECT  3.720 0.830 3.840 1.140 ;
        RECT  3.700 0.310 3.790 0.690 ;
        RECT  3.610 0.830 3.720 0.940 ;
        RECT  3.590 0.310 3.700 0.420 ;
        RECT  3.520 0.530 3.610 0.940 ;
        RECT  3.430 0.275 3.500 0.385 ;
        RECT  3.430 1.035 3.490 1.165 ;
        RECT  3.350 1.255 3.440 1.505 ;
        RECT  3.340 0.275 3.430 1.165 ;
        RECT  1.340 1.255 3.350 1.345 ;
        RECT  3.330 0.275 3.340 0.595 ;
        RECT  2.895 0.995 3.340 1.165 ;
        RECT  2.740 0.725 3.250 0.895 ;
        RECT  2.595 0.305 2.740 1.145 ;
        RECT  2.540 1.035 2.595 1.145 ;
        RECT  1.035 0.275 2.485 0.385 ;
        RECT  1.085 1.435 2.445 1.525 ;
        RECT  2.260 0.510 2.360 1.145 ;
        RECT  2.045 0.510 2.260 0.645 ;
        RECT  2.035 1.025 2.260 1.145 ;
        RECT  1.945 0.750 2.030 0.920 ;
        RECT  1.855 0.490 1.945 1.145 ;
        RECT  1.550 0.490 1.855 0.600 ;
        RECT  1.520 1.030 1.855 1.145 ;
        RECT  1.235 0.900 1.340 1.345 ;
        RECT  1.010 0.685 1.100 1.305 ;
        RECT  0.830 1.395 1.085 1.525 ;
        RECT  0.920 0.275 1.035 0.525 ;
        RECT  0.190 1.215 1.010 1.305 ;
        RECT  0.705 0.475 0.810 1.125 ;
        RECT  0.650 0.475 0.705 0.665 ;
        RECT  0.555 1.010 0.705 1.125 ;
        RECT  0.155 0.285 0.195 0.460 ;
        RECT  0.155 1.215 0.190 1.515 ;
        RECT  0.045 0.285 0.155 1.515 ;
    END
END EDFQD4

MACRO FA1D0
    CLASS CORE ;
    FOREIGN FA1D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.510 4.550 1.155 ;
        RECT  4.400 0.510 4.450 0.620 ;
        RECT  4.400 1.045 4.450 1.155 ;
        RECT  4.290 0.275 4.400 0.620 ;
        RECT  4.300 1.045 4.400 1.255 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.825 0.275 4.950 1.290 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.0529 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.510 3.965 0.890 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0928 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.580 0.710 1.650 0.940 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 -0.165 5.000 0.165 ;
        RECT  4.515 -0.165 4.700 0.420 ;
        RECT  0.475 -0.165 4.515 0.165 ;
        RECT  0.305 -0.165 0.475 0.400 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.825 1.635 5.000 1.965 ;
        RECT  1.655 1.440 1.825 1.965 ;
        RECT  0.475 1.635 1.655 1.965 ;
        RECT  0.305 1.390 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.640 0.730 4.735 1.515 ;
        RECT  2.605 1.425 4.640 1.515 ;
        RECT  4.210 0.775 4.360 0.895 ;
        RECT  4.120 0.775 4.210 1.335 ;
        RECT  3.740 0.310 4.190 0.420 ;
        RECT  3.180 1.245 4.120 1.335 ;
        RECT  3.740 0.985 4.030 1.155 ;
        RECT  3.650 0.275 3.740 1.155 ;
        RECT  2.980 0.275 3.650 0.365 ;
        RECT  3.540 0.730 3.650 0.940 ;
        RECT  3.450 0.475 3.560 0.585 ;
        RECT  3.360 0.475 3.450 1.155 ;
        RECT  3.280 1.045 3.360 1.155 ;
        RECT  3.180 0.475 3.250 0.665 ;
        RECT  3.090 0.475 3.180 1.335 ;
        RECT  2.975 1.205 3.090 1.335 ;
        RECT  2.870 0.275 2.980 0.880 ;
        RECT  2.865 0.790 2.870 0.880 ;
        RECT  2.755 0.790 2.865 1.335 ;
        RECT  2.610 0.275 2.720 0.615 ;
        RECT  2.605 0.505 2.610 0.615 ;
        RECT  2.495 0.505 2.605 1.515 ;
        RECT  2.290 0.455 2.390 1.350 ;
        RECT  1.510 1.240 2.290 1.350 ;
        RECT  2.080 0.275 2.180 1.150 ;
        RECT  2.025 0.275 2.080 0.675 ;
        RECT  1.920 1.040 2.080 1.150 ;
        RECT  1.840 0.275 1.935 0.930 ;
        RECT  0.990 0.275 1.840 0.365 ;
        RECT  1.470 0.455 1.585 0.565 ;
        RECT  1.470 1.040 1.510 1.470 ;
        RECT  1.380 0.455 1.470 1.470 ;
        RECT  1.320 0.775 1.380 0.945 ;
        RECT  1.210 0.455 1.270 0.625 ;
        RECT  1.210 1.055 1.255 1.525 ;
        RECT  1.120 0.455 1.210 1.525 ;
        RECT  0.710 1.435 1.120 1.525 ;
        RECT  0.880 0.275 0.990 1.325 ;
        RECT  0.705 0.580 0.755 1.120 ;
        RECT  0.620 1.210 0.710 1.525 ;
        RECT  0.645 0.270 0.705 1.120 ;
        RECT  0.595 0.270 0.645 0.690 ;
        RECT  0.545 1.015 0.645 1.120 ;
        RECT  0.360 1.210 0.620 1.300 ;
        RECT  0.360 0.755 0.520 0.925 ;
        RECT  0.270 0.490 0.360 1.300 ;
        RECT  0.185 0.490 0.270 0.590 ;
        RECT  0.185 1.210 0.270 1.300 ;
        RECT  0.075 0.370 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.420 ;
    END
END FA1D0

MACRO FA1D1
    CLASS CORE ;
    FOREIGN FA1D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1390 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.045 0.300 5.155 1.190 ;
        RECT  4.890 0.485 5.045 0.615 ;
        RECT  4.855 1.080 5.045 1.190 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.445 0.285 5.550 1.510 ;
        RECT  5.425 0.285 5.445 0.675 ;
        RECT  5.425 1.050 5.445 1.510 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.645 0.280 4.765 0.695 ;
        RECT  4.555 0.585 4.645 0.695 ;
        RECT  4.445 0.585 4.555 0.905 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0914 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.710 1.355 0.925 ;
        RECT  1.050 0.480 1.160 0.925 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.440 0.895 ;
        RECT  0.050 0.690 0.150 1.110 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 5.600 0.165 ;
        RECT  0.075 -0.165 0.185 0.475 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.635 5.600 1.965 ;
        RECT  5.100 1.500 5.270 1.965 ;
        RECT  0.185 1.635 5.100 1.965 ;
        RECT  0.075 1.305 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.245 0.725 5.335 1.390 ;
        RECT  4.990 1.300 5.245 1.390 ;
        RECT  4.890 1.300 4.990 1.505 ;
        RECT  4.765 0.825 4.945 0.935 ;
        RECT  3.135 1.415 4.890 1.505 ;
        RECT  4.675 0.825 4.765 1.325 ;
        RECT  3.695 1.235 4.675 1.325 ;
        RECT  4.440 0.275 4.550 0.495 ;
        RECT  4.245 1.015 4.525 1.125 ;
        RECT  4.245 0.275 4.440 0.365 ;
        RECT  4.155 0.275 4.245 1.125 ;
        RECT  3.495 0.275 4.155 0.365 ;
        RECT  4.025 0.735 4.155 0.905 ;
        RECT  3.935 0.475 4.065 0.600 ;
        RECT  3.935 1.015 4.005 1.125 ;
        RECT  3.845 0.475 3.935 1.125 ;
        RECT  3.795 1.015 3.845 1.125 ;
        RECT  3.695 0.460 3.755 0.875 ;
        RECT  3.645 0.460 3.695 1.325 ;
        RECT  3.585 0.765 3.645 1.325 ;
        RECT  3.500 1.195 3.585 1.325 ;
        RECT  3.400 0.275 3.495 0.910 ;
        RECT  3.395 0.275 3.400 1.305 ;
        RECT  3.290 0.810 3.395 1.305 ;
        RECT  3.145 0.330 3.255 0.660 ;
        RECT  3.135 0.550 3.145 0.660 ;
        RECT  3.040 0.550 3.135 1.505 ;
        RECT  2.750 0.275 3.040 0.415 ;
        RECT  2.860 0.525 2.950 1.485 ;
        RECT  2.225 1.375 2.860 1.485 ;
        RECT  2.660 0.275 2.750 1.190 ;
        RECT  2.620 0.275 2.660 0.415 ;
        RECT  2.505 1.080 2.660 1.190 ;
        RECT  2.480 0.530 2.570 0.945 ;
        RECT  2.460 0.275 2.480 0.945 ;
        RECT  2.370 0.275 2.460 0.640 ;
        RECT  1.680 0.275 2.370 0.365 ;
        RECT  2.115 0.475 2.225 1.485 ;
        RECT  1.970 0.755 2.115 0.925 ;
        RECT  2.000 1.375 2.115 1.485 ;
        RECT  1.880 0.475 1.975 0.645 ;
        RECT  1.885 1.035 1.940 1.205 ;
        RECT  1.880 1.035 1.885 1.525 ;
        RECT  1.790 0.475 1.880 1.525 ;
        RECT  0.650 1.435 1.790 1.525 ;
        RECT  1.570 0.275 1.680 1.325 ;
        RECT  1.270 0.285 1.450 0.600 ;
        RECT  0.960 1.135 1.450 1.245 ;
        RECT  0.960 0.285 1.270 0.375 ;
        RECT  0.870 0.285 0.960 1.245 ;
        RECT  0.830 0.285 0.870 0.675 ;
        RECT  0.790 1.085 0.870 1.245 ;
        RECT  0.650 0.775 0.780 0.945 ;
        RECT  0.560 0.575 0.650 1.525 ;
        RECT  0.445 0.575 0.560 0.675 ;
        RECT  0.445 1.025 0.560 1.135 ;
        RECT  0.335 0.285 0.445 0.675 ;
        RECT  0.335 1.025 0.445 1.525 ;
    END
END FA1D1

MACRO FA1D2
    CLASS CORE ;
    FOREIGN FA1D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.965 0.545 5.065 1.290 ;
        RECT  4.835 0.285 4.965 0.675 ;
        RECT  4.835 1.110 4.965 1.290 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.510 5.555 1.495 ;
        RECT  5.445 0.275 5.475 1.495 ;
        RECT  5.365 0.275 5.445 0.675 ;
        RECT  5.365 1.055 5.445 1.495 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.510 4.555 0.905 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.710 1.355 0.925 ;
        RECT  1.050 0.480 1.160 0.925 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.430 0.895 ;
        RECT  0.050 0.690 0.150 1.110 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.255 0.810 5.355 0.910 ;
        RECT  5.155 0.810 5.255 1.515 ;
        RECT  3.130 1.415 5.155 1.515 ;
        RECT  4.745 0.805 4.870 0.915 ;
        RECT  4.645 0.805 4.745 1.325 ;
        RECT  3.685 1.235 4.645 1.325 ;
        RECT  4.235 0.275 4.515 0.420 ;
        RECT  4.235 1.015 4.515 1.125 ;
        RECT  4.145 0.275 4.235 1.125 ;
        RECT  3.440 0.275 4.145 0.365 ;
        RECT  4.015 0.735 4.145 0.905 ;
        RECT  3.925 0.475 4.015 0.600 ;
        RECT  3.925 1.015 3.995 1.125 ;
        RECT  3.835 0.475 3.925 1.125 ;
        RECT  3.785 1.015 3.835 1.125 ;
        RECT  3.685 0.455 3.700 0.905 ;
        RECT  3.590 0.455 3.685 1.325 ;
        RECT  3.575 0.805 3.590 1.325 ;
        RECT  3.510 1.195 3.575 1.325 ;
        RECT  3.390 0.275 3.440 0.905 ;
        RECT  3.390 1.200 3.420 1.325 ;
        RECT  3.340 0.275 3.390 1.325 ;
        RECT  3.280 0.805 3.340 1.325 ;
        RECT  3.240 1.200 3.280 1.325 ;
        RECT  3.145 0.545 3.230 0.655 ;
        RECT  3.130 0.545 3.145 0.905 ;
        RECT  3.050 0.545 3.130 1.515 ;
        RECT  3.030 0.805 3.050 1.515 ;
        RECT  2.740 0.275 3.025 0.415 ;
        RECT  2.830 0.505 2.940 1.485 ;
        RECT  2.215 1.375 2.830 1.485 ;
        RECT  2.650 0.275 2.740 1.190 ;
        RECT  2.600 0.275 2.650 0.415 ;
        RECT  2.505 1.080 2.650 1.190 ;
        RECT  2.470 0.735 2.560 0.945 ;
        RECT  2.360 0.275 2.470 0.945 ;
        RECT  1.670 0.275 2.360 0.365 ;
        RECT  2.105 0.475 2.215 1.485 ;
        RECT  1.960 0.755 2.105 0.925 ;
        RECT  1.990 1.375 2.105 1.485 ;
        RECT  1.870 0.475 1.985 0.645 ;
        RECT  1.875 1.035 1.960 1.205 ;
        RECT  1.870 1.035 1.875 1.525 ;
        RECT  1.780 0.475 1.870 1.525 ;
        RECT  0.435 1.435 1.780 1.525 ;
        RECT  1.560 0.275 1.670 1.325 ;
        RECT  1.260 0.285 1.440 0.600 ;
        RECT  0.950 1.135 1.440 1.245 ;
        RECT  0.950 0.285 1.260 0.375 ;
        RECT  0.860 0.285 0.950 1.245 ;
        RECT  0.820 0.285 0.860 0.675 ;
        RECT  0.780 1.085 0.860 1.245 ;
        RECT  0.640 0.775 0.770 0.945 ;
        RECT  0.550 0.575 0.640 1.135 ;
        RECT  0.435 0.575 0.550 0.675 ;
        RECT  0.435 1.025 0.550 1.135 ;
        RECT  0.325 0.285 0.435 0.675 ;
        RECT  0.325 1.025 0.435 1.525 ;
    END
END FA1D2

MACRO FA1D4
    CLASS CORE ;
    FOREIGN FA1D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 1.100 6.635 1.300 ;
        RECT  6.450 0.300 6.625 0.500 ;
        RECT  6.150 0.300 6.450 1.300 ;
        RECT  6.015 0.300 6.150 0.500 ;
        RECT  6.020 1.100 6.150 1.300 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.555 0.265 7.665 0.680 ;
        RECT  7.555 1.040 7.665 1.470 ;
        RECT  7.450 0.570 7.555 0.680 ;
        RECT  7.450 1.040 7.555 1.150 ;
        RECT  7.150 0.570 7.450 1.150 ;
        RECT  7.145 0.570 7.150 0.680 ;
        RECT  7.145 1.040 7.150 1.150 ;
        RECT  7.035 0.265 7.145 0.680 ;
        RECT  7.035 1.040 7.145 1.470 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.1101 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.700 5.750 0.900 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.1437 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.950 1.100 ;
        RECT  2.805 0.710 2.850 0.925 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.350 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.925 -0.165 8.000 0.165 ;
        RECT  7.815 -0.165 7.925 0.695 ;
        RECT  7.405 -0.165 7.815 0.165 ;
        RECT  7.295 -0.165 7.405 0.480 ;
        RECT  6.885 -0.165 7.295 0.165 ;
        RECT  6.775 -0.165 6.885 0.665 ;
        RECT  5.865 -0.165 6.775 0.165 ;
        RECT  5.755 -0.165 5.865 0.505 ;
        RECT  0.000 -0.165 5.755 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.925 1.635 8.000 1.965 ;
        RECT  7.815 1.040 7.925 1.965 ;
        RECT  7.405 1.635 7.815 1.965 ;
        RECT  7.295 1.260 7.405 1.965 ;
        RECT  0.000 1.635 7.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.555 0.265 7.665 0.680 ;
        RECT  7.555 1.040 7.665 1.470 ;
        RECT  7.550 0.570 7.555 0.680 ;
        RECT  7.550 1.040 7.555 1.150 ;
        RECT  7.035 0.265 7.050 0.680 ;
        RECT  7.035 1.040 7.050 1.470 ;
        RECT  6.550 1.100 6.635 1.300 ;
        RECT  6.550 0.300 6.625 0.500 ;
        RECT  6.015 0.300 6.050 0.500 ;
        RECT  6.020 1.100 6.050 1.300 ;
        RECT  6.880 0.780 7.040 0.890 ;
        RECT  6.790 0.780 6.880 1.495 ;
        RECT  3.790 1.405 6.790 1.495 ;
        RECT  5.930 0.780 6.030 0.890 ;
        RECT  5.840 0.780 5.930 1.315 ;
        RECT  4.320 1.225 5.840 1.315 ;
        RECT  5.360 0.455 5.655 0.565 ;
        RECT  5.360 1.025 5.655 1.135 ;
        RECT  5.265 0.275 5.360 1.135 ;
        RECT  4.110 0.275 5.265 0.365 ;
        RECT  4.920 0.765 5.265 0.875 ;
        RECT  4.570 0.485 5.155 0.595 ;
        RECT  4.570 1.025 5.115 1.135 ;
        RECT  4.480 0.485 4.570 1.135 ;
        RECT  4.410 1.025 4.480 1.135 ;
        RECT  4.320 0.455 4.370 0.625 ;
        RECT  4.230 0.455 4.320 1.315 ;
        RECT  4.110 1.190 4.230 1.315 ;
        RECT  4.010 0.275 4.110 0.880 ;
        RECT  4.000 0.275 4.010 1.315 ;
        RECT  3.900 0.790 4.000 1.315 ;
        RECT  3.790 0.495 3.900 0.605 ;
        RECT  3.700 0.495 3.790 1.495 ;
        RECT  3.650 1.210 3.700 1.495 ;
        RECT  3.540 0.465 3.590 0.645 ;
        RECT  3.490 0.465 3.540 1.340 ;
        RECT  2.205 0.275 3.500 0.375 ;
        RECT  3.450 0.465 3.490 1.530 ;
        RECT  3.380 1.250 3.450 1.530 ;
        RECT  2.725 1.250 3.380 1.340 ;
        RECT  3.250 0.520 3.360 1.135 ;
        RECT  3.085 0.520 3.250 0.630 ;
        RECT  3.090 1.025 3.250 1.135 ;
        RECT  2.700 0.485 2.800 0.595 ;
        RECT  2.700 1.035 2.725 1.465 ;
        RECT  2.610 0.485 2.700 1.465 ;
        RECT  2.520 0.775 2.610 0.945 ;
        RECT  2.420 0.485 2.520 0.595 ;
        RECT  2.420 1.060 2.470 1.525 ;
        RECT  2.330 0.485 2.420 1.525 ;
        RECT  0.685 1.435 2.330 1.525 ;
        RECT  2.095 0.275 2.205 1.330 ;
        RECT  1.415 1.235 1.985 1.345 ;
        RECT  1.835 0.275 1.945 0.550 ;
        RECT  1.685 0.785 1.870 0.895 ;
        RECT  1.415 0.275 1.835 0.365 ;
        RECT  1.675 1.035 1.735 1.145 ;
        RECT  1.675 0.455 1.685 0.895 ;
        RECT  1.575 0.455 1.675 1.145 ;
        RECT  1.525 1.035 1.575 1.145 ;
        RECT  1.325 0.275 1.415 1.345 ;
        RECT  1.025 0.485 1.325 0.595 ;
        RECT  1.025 1.235 1.325 1.345 ;
        RECT  0.685 0.780 1.235 0.895 ;
        RECT  0.575 0.275 0.685 1.525 ;
        RECT  0.185 0.465 0.575 0.575 ;
        RECT  0.185 1.025 0.575 1.115 ;
        RECT  0.075 0.365 0.185 0.575 ;
        RECT  0.075 1.025 0.185 1.470 ;
    END
END FA1D4

MACRO FCICIND1
    CLASS CORE ;
    FOREIGN FCICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CO
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.555 2.155 1.290 ;
        RECT  1.965 0.555 2.045 0.690 ;
        RECT  1.820 1.110 2.045 1.290 ;
        RECT  1.845 0.275 1.965 0.690 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.710 2.370 1.100 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.0857 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.635 1.235 0.965 ;
        RECT  0.750 0.635 1.125 0.725 ;
        RECT  0.645 0.635 0.750 1.090 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0993 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.550 1.090 ;
        RECT  0.290 0.815 0.450 1.005 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 -0.165 2.600 0.165 ;
        RECT  2.140 -0.165 2.250 0.445 ;
        RECT  0.840 -0.165 2.140 0.165 ;
        RECT  0.670 -0.165 0.840 0.365 ;
        RECT  0.000 -0.165 0.670 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.635 2.600 1.965 ;
        RECT  0.625 1.200 0.750 1.965 ;
        RECT  0.000 1.635 0.625 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.460 0.325 2.550 1.525 ;
        RECT  2.425 0.325 2.460 0.585 ;
        RECT  2.405 1.235 2.460 1.525 ;
        RECT  0.950 1.435 2.405 1.525 ;
        RECT  1.435 0.800 1.935 0.910 ;
        RECT  1.565 0.275 1.695 0.570 ;
        RECT  1.580 1.090 1.680 1.345 ;
        RECT  1.160 1.255 1.580 1.345 ;
        RECT  0.980 0.275 1.565 0.365 ;
        RECT  1.435 1.075 1.470 1.165 ;
        RECT  1.325 0.455 1.435 1.165 ;
        RECT  0.200 0.455 1.325 0.545 ;
        RECT  1.270 1.075 1.325 1.165 ;
        RECT  1.060 1.090 1.160 1.345 ;
        RECT  0.950 0.815 1.005 1.005 ;
        RECT  0.860 0.815 0.950 1.525 ;
        RECT  0.065 0.325 0.200 1.515 ;
    END
END FCICIND1

MACRO FCICIND2
    CLASS CORE ;
    FOREIGN FCICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CO
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.580 2.355 1.300 ;
        RECT  2.165 0.580 2.245 0.690 ;
        RECT  2.010 1.110 2.245 1.300 ;
        RECT  2.045 0.275 2.165 0.690 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.710 2.570 1.100 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.0857 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.635 1.235 0.965 ;
        RECT  0.750 0.635 1.125 0.725 ;
        RECT  0.645 0.635 0.750 1.090 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0993 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.550 1.090 ;
        RECT  0.290 0.815 0.450 1.005 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 -0.165 2.800 0.165 ;
        RECT  2.340 -0.165 2.450 0.465 ;
        RECT  0.840 -0.165 2.340 0.165 ;
        RECT  0.670 -0.165 0.840 0.365 ;
        RECT  0.000 -0.165 0.670 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.635 2.800 1.965 ;
        RECT  0.645 1.200 0.750 1.965 ;
        RECT  0.000 1.635 0.645 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.660 0.325 2.750 1.525 ;
        RECT  2.625 0.325 2.660 0.580 ;
        RECT  2.605 1.235 2.660 1.525 ;
        RECT  0.950 1.435 2.605 1.525 ;
        RECT  1.435 0.785 2.135 0.895 ;
        RECT  1.565 0.275 1.695 0.580 ;
        RECT  1.580 1.080 1.695 1.345 ;
        RECT  1.160 1.255 1.580 1.345 ;
        RECT  0.980 0.275 1.565 0.365 ;
        RECT  1.435 1.075 1.470 1.165 ;
        RECT  1.325 0.455 1.435 1.165 ;
        RECT  0.200 0.455 1.325 0.545 ;
        RECT  1.270 1.075 1.325 1.165 ;
        RECT  1.060 1.080 1.160 1.345 ;
        RECT  0.950 0.815 1.005 1.005 ;
        RECT  0.860 0.815 0.950 1.525 ;
        RECT  0.065 0.325 0.200 1.515 ;
    END
END FCICIND2

MACRO FCICOND1
    CLASS CORE ;
    FOREIGN FCICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CON
        ANTENNADIFFAREA 0.3110 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.455 1.355 1.290 ;
        RECT  0.195 0.455 1.245 0.545 ;
        RECT  0.150 0.310 0.195 0.545 ;
        RECT  0.150 1.200 0.175 1.490 ;
        RECT  0.050 0.310 0.150 1.490 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.955 1.090 ;
        RECT  0.740 0.710 0.845 0.945 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0891 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.655 1.155 1.290 ;
        RECT  0.555 1.200 1.045 1.290 ;
        RECT  0.555 0.710 0.620 0.945 ;
        RECT  0.445 0.710 0.555 1.290 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1077 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.655 0.355 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.165 1.800 0.165 ;
        RECT  0.590 -0.165 0.760 0.365 ;
        RECT  0.000 -0.165 0.590 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.635 1.800 1.965 ;
        RECT  0.590 1.395 0.780 1.965 ;
        RECT  0.000 1.635 0.590 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.495 0.275 1.605 0.685 ;
        RECT  1.495 1.015 1.605 1.510 ;
        RECT  0.900 0.275 1.495 0.365 ;
        RECT  0.900 1.400 1.495 1.510 ;
    END
END FCICOND1

MACRO FCICOND2
    CLASS CORE ;
    FOREIGN FCICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CON
        ANTENNADIFFAREA 0.1860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.465 0.545 2.555 1.195 ;
        RECT  2.445 0.275 2.465 1.505 ;
        RECT  2.355 0.275 2.445 0.675 ;
        RECT  2.355 1.055 2.445 1.505 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.955 1.090 ;
        RECT  0.740 0.710 0.845 0.945 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0891 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.655 1.155 1.290 ;
        RECT  0.555 1.200 1.045 1.290 ;
        RECT  0.555 0.710 0.620 0.945 ;
        RECT  0.445 0.710 0.555 1.290 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1077 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.655 0.355 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.725 -0.165 2.800 0.165 ;
        RECT  2.615 -0.165 2.725 0.455 ;
        RECT  2.170 -0.165 2.615 0.165 ;
        RECT  2.060 -0.165 2.170 0.675 ;
        RECT  0.760 -0.165 2.060 0.165 ;
        RECT  0.590 -0.165 0.760 0.365 ;
        RECT  0.000 -0.165 0.590 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.725 1.635 2.800 1.965 ;
        RECT  2.615 1.285 2.725 1.965 ;
        RECT  2.165 1.635 2.615 1.965 ;
        RECT  2.055 1.055 2.165 1.965 ;
        RECT  0.780 1.635 2.055 1.965 ;
        RECT  0.590 1.395 0.780 1.965 ;
        RECT  0.000 1.635 0.590 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.950 0.765 2.275 0.935 ;
        RECT  1.865 0.535 1.950 1.195 ;
        RECT  1.850 0.275 1.865 1.490 ;
        RECT  1.755 0.275 1.850 0.685 ;
        RECT  1.355 0.800 1.760 0.900 ;
        RECT  1.495 0.275 1.605 0.685 ;
        RECT  1.495 1.015 1.605 1.500 ;
        RECT  0.900 0.275 1.495 0.365 ;
        RECT  0.900 1.380 1.495 1.500 ;
        RECT  1.245 0.455 1.355 1.270 ;
        RECT  0.195 0.455 1.245 0.545 ;
        RECT  0.150 0.310 0.195 0.545 ;
        RECT  0.150 1.200 0.175 1.490 ;
        RECT  0.050 0.310 0.150 1.490 ;
        RECT  1.755 1.015 1.850 1.490 ;
    END
END FCICOND2

MACRO FCSICIND1
    CLASS CORE ;
    FOREIGN FCSICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.850 0.310 9.950 1.490 ;
        RECT  9.815 0.310 9.850 0.575 ;
        RECT  9.820 1.040 9.850 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0921 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.440 0.700 9.550 1.100 ;
        RECT  9.410 0.700 9.440 0.940 ;
        END
    END CS
    PIN CO1
        ANTENNADIFFAREA 0.1490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.550 0.635 5.690 0.725 ;
        RECT  5.550 1.120 5.610 1.290 ;
        RECT  5.450 0.635 5.550 1.290 ;
        END
    END CO1
    PIN CO0
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.635 5.350 1.290 ;
        RECT  5.110 0.635 5.250 0.725 ;
        RECT  5.195 1.120 5.250 1.290 ;
        END
    END CO0
    PIN CIN1
        ANTENNAGATEAREA 0.0529 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.440 0.710 7.780 0.890 ;
        END
    END CIN1
    PIN CIN0
        ANTENNAGATEAREA 0.0530 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CIN0
    PIN B
        ANTENNAGATEAREA 0.0927 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.350 1.100 ;
        RECT  1.195 0.700 1.250 0.940 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.430 0.895 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.650 -0.165 10.000 0.165 ;
        RECT  9.505 -0.165 9.650 0.575 ;
        RECT  0.000 -0.165 9.505 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 10.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.730 0.730 9.760 0.920 ;
        RECT  9.640 0.730 9.730 1.525 ;
        RECT  8.785 1.435 9.640 1.525 ;
        RECT  9.260 0.310 9.360 0.575 ;
        RECT  9.260 1.035 9.345 1.335 ;
        RECT  9.235 0.310 9.260 1.335 ;
        RECT  9.160 0.465 9.235 1.125 ;
        RECT  8.985 1.235 9.095 1.345 ;
        RECT  8.985 0.275 9.070 0.865 ;
        RECT  8.970 0.275 8.985 1.345 ;
        RECT  3.590 0.275 8.970 0.365 ;
        RECT  8.895 0.775 8.970 1.345 ;
        RECT  8.785 0.520 8.870 0.630 ;
        RECT  8.675 0.520 8.785 1.525 ;
        RECT  8.500 1.180 8.525 1.495 ;
        RECT  8.385 0.455 8.500 1.495 ;
        RECT  7.070 1.385 8.385 1.495 ;
        RECT  8.205 0.455 8.295 1.295 ;
        RECT  8.120 0.455 8.205 0.640 ;
        RECT  6.945 1.205 8.205 1.295 ;
        RECT  8.020 0.750 8.095 0.920 ;
        RECT  7.930 0.490 8.020 1.115 ;
        RECT  7.555 0.490 7.930 0.600 ;
        RECT  7.405 1.015 7.930 1.115 ;
        RECT  7.285 0.490 7.450 0.600 ;
        RECT  7.195 0.490 7.285 1.115 ;
        RECT  7.070 1.015 7.195 1.115 ;
        RECT  6.995 0.455 7.105 0.875 ;
        RECT  6.945 0.785 6.995 0.875 ;
        RECT  6.845 0.785 6.945 1.295 ;
        RECT  6.755 0.495 6.885 0.605 ;
        RECT  6.665 0.495 6.755 1.295 ;
        RECT  5.810 1.205 6.665 1.295 ;
        RECT  6.465 0.475 6.575 1.115 ;
        RECT  6.265 1.385 6.475 1.500 ;
        RECT  6.260 1.005 6.465 1.115 ;
        RECT  6.270 0.675 6.340 0.885 ;
        RECT  6.170 0.460 6.270 0.885 ;
        RECT  4.540 1.400 6.265 1.500 ;
        RECT  6.160 0.460 6.170 1.115 ;
        RECT  6.080 0.785 6.160 1.115 ;
        RECT  5.980 1.025 6.080 1.115 ;
        RECT  5.900 0.455 5.990 0.915 ;
        RECT  4.905 0.455 5.900 0.545 ;
        RECT  5.720 0.845 5.810 1.295 ;
        RECT  5.650 0.845 5.720 1.015 ;
        RECT  5.085 0.845 5.160 1.015 ;
        RECT  4.995 0.845 5.085 1.295 ;
        RECT  4.150 1.205 4.995 1.295 ;
        RECT  4.815 0.455 4.905 0.915 ;
        RECT  4.725 1.025 4.825 1.115 ;
        RECT  4.650 0.785 4.725 1.115 ;
        RECT  4.635 0.475 4.650 1.115 ;
        RECT  4.475 0.475 4.635 0.895 ;
        RECT  4.350 1.005 4.545 1.115 ;
        RECT  4.330 1.385 4.540 1.500 ;
        RECT  4.240 0.475 4.350 1.115 ;
        RECT  2.190 1.400 4.330 1.500 ;
        RECT  4.060 0.665 4.150 1.295 ;
        RECT  4.040 0.665 4.060 0.755 ;
        RECT  3.930 0.465 4.040 0.755 ;
        RECT  3.860 0.845 3.960 1.295 ;
        RECT  3.790 0.845 3.860 0.935 ;
        RECT  2.495 1.205 3.860 1.295 ;
        RECT  3.680 0.455 3.790 0.935 ;
        RECT  3.590 1.025 3.735 1.115 ;
        RECT  3.500 0.275 3.590 1.115 ;
        RECT  3.365 0.490 3.500 0.600 ;
        RECT  1.670 0.275 3.410 0.385 ;
        RECT  2.940 1.015 3.390 1.115 ;
        RECT  2.940 0.490 3.275 0.600 ;
        RECT  2.850 0.490 2.940 1.115 ;
        RECT  2.630 0.780 2.850 0.890 ;
        RECT  2.495 0.535 2.740 0.645 ;
        RECT  2.405 0.535 2.495 1.295 ;
        RECT  2.190 0.535 2.265 0.645 ;
        RECT  2.080 0.535 2.190 1.500 ;
        RECT  2.075 0.535 2.080 0.945 ;
        RECT  2.000 0.775 2.075 0.945 ;
        RECT  1.890 0.535 1.985 0.645 ;
        RECT  1.890 1.045 1.935 1.525 ;
        RECT  1.800 0.535 1.890 1.525 ;
        RECT  0.670 1.435 1.800 1.525 ;
        RECT  1.560 0.275 1.670 1.330 ;
        RECT  1.080 1.235 1.450 1.345 ;
        RECT  1.300 0.340 1.410 0.590 ;
        RECT  1.080 0.500 1.300 0.590 ;
        RECT  0.990 0.500 1.080 1.345 ;
        RECT  0.935 0.500 0.990 0.675 ;
        RECT  0.780 1.235 0.990 1.345 ;
        RECT  0.820 0.265 0.935 0.675 ;
        RECT  0.670 0.780 0.880 0.895 ;
        RECT  0.580 0.575 0.670 1.525 ;
        RECT  0.445 0.575 0.580 0.675 ;
        RECT  0.445 1.425 0.580 1.525 ;
        RECT  0.315 0.265 0.445 0.675 ;
        RECT  0.315 1.040 0.445 1.525 ;
    END
END FCSICIND1

MACRO FCSICIND2
    CLASS CORE ;
    FOREIGN FCSICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.050 0.310 10.150 1.490 ;
        RECT  10.015 0.310 10.050 0.520 ;
        RECT  10.020 1.040 10.050 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0925 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.650 0.700 9.750 1.100 ;
        RECT  9.620 0.700 9.650 0.940 ;
        END
    END CS
    PIN CO1
        ANTENNADIFFAREA 0.1800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.755 0.635 5.935 0.725 ;
        RECT  5.755 1.120 5.865 1.295 ;
        RECT  5.650 0.635 5.755 1.295 ;
        END
    END CO1
    PIN CO0
        ANTENNADIFFAREA 0.1800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.635 5.350 1.295 ;
        RECT  5.125 0.635 5.250 0.725 ;
        RECT  5.195 1.120 5.250 1.295 ;
        END
    END CO0
    PIN CIN1
        ANTENNAGATEAREA 0.0527 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.710 8.035 0.890 ;
        END
    END CIN1
    PIN CIN0
        ANTENNAGATEAREA 0.0530 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CIN0
    PIN B
        ANTENNAGATEAREA 0.0927 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.350 1.100 ;
        RECT  1.195 0.700 1.250 0.940 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.430 0.895 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.845 -0.165 10.200 0.165 ;
        RECT  9.745 -0.165 9.845 0.575 ;
        RECT  0.000 -0.165 9.745 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 10.200 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.930 0.730 9.960 0.940 ;
        RECT  9.840 0.730 9.930 1.525 ;
        RECT  8.995 1.435 9.840 1.525 ;
        RECT  9.480 0.415 9.625 0.525 ;
        RECT  9.480 1.035 9.560 1.335 ;
        RECT  9.455 0.415 9.480 1.335 ;
        RECT  9.370 0.415 9.455 1.125 ;
        RECT  9.180 0.275 9.280 1.345 ;
        RECT  3.590 0.275 9.180 0.365 ;
        RECT  9.140 1.115 9.180 1.345 ;
        RECT  8.995 0.520 9.080 0.630 ;
        RECT  8.885 0.520 8.995 1.525 ;
        RECT  8.710 1.180 8.735 1.495 ;
        RECT  8.595 0.455 8.710 1.495 ;
        RECT  7.325 1.385 8.595 1.495 ;
        RECT  8.415 0.455 8.505 1.295 ;
        RECT  8.330 0.455 8.415 0.640 ;
        RECT  7.200 1.205 8.415 1.295 ;
        RECT  8.240 0.750 8.305 0.920 ;
        RECT  8.145 0.490 8.240 1.115 ;
        RECT  7.790 0.490 8.145 0.600 ;
        RECT  7.650 1.015 8.145 1.115 ;
        RECT  7.540 0.490 7.680 0.600 ;
        RECT  7.450 0.490 7.540 1.115 ;
        RECT  7.325 1.015 7.450 1.115 ;
        RECT  7.250 0.455 7.360 0.875 ;
        RECT  7.200 0.785 7.250 0.875 ;
        RECT  7.100 0.785 7.200 1.295 ;
        RECT  7.010 0.495 7.140 0.605 ;
        RECT  6.920 0.495 7.010 1.295 ;
        RECT  6.065 1.205 6.920 1.295 ;
        RECT  6.720 0.475 6.830 1.115 ;
        RECT  2.190 1.385 6.730 1.485 ;
        RECT  6.515 1.005 6.720 1.115 ;
        RECT  6.525 0.675 6.595 0.885 ;
        RECT  6.425 0.460 6.525 0.885 ;
        RECT  6.415 0.460 6.425 1.115 ;
        RECT  6.335 0.785 6.415 1.115 ;
        RECT  6.235 1.025 6.335 1.115 ;
        RECT  6.155 0.455 6.245 0.915 ;
        RECT  4.905 0.455 6.155 0.545 ;
        RECT  5.975 0.845 6.065 1.295 ;
        RECT  5.905 0.845 5.975 1.015 ;
        RECT  5.085 0.845 5.160 1.015 ;
        RECT  4.995 0.845 5.085 1.295 ;
        RECT  4.150 1.205 4.995 1.295 ;
        RECT  4.815 0.455 4.905 0.915 ;
        RECT  4.725 1.025 4.825 1.115 ;
        RECT  4.650 0.785 4.725 1.115 ;
        RECT  4.635 0.475 4.650 1.115 ;
        RECT  4.475 0.475 4.635 0.895 ;
        RECT  4.350 1.005 4.545 1.115 ;
        RECT  4.240 0.475 4.350 1.115 ;
        RECT  4.060 0.665 4.150 1.295 ;
        RECT  4.040 0.665 4.060 0.755 ;
        RECT  3.930 0.465 4.040 0.755 ;
        RECT  3.860 0.845 3.960 1.295 ;
        RECT  3.790 0.845 3.860 0.935 ;
        RECT  2.495 1.205 3.860 1.295 ;
        RECT  3.680 0.455 3.790 0.935 ;
        RECT  3.590 1.025 3.735 1.115 ;
        RECT  3.500 0.275 3.590 1.115 ;
        RECT  3.365 0.490 3.500 0.600 ;
        RECT  1.670 0.275 3.410 0.385 ;
        RECT  2.940 1.015 3.390 1.115 ;
        RECT  2.940 0.490 3.275 0.600 ;
        RECT  2.850 0.490 2.940 1.115 ;
        RECT  2.630 0.780 2.850 0.890 ;
        RECT  2.495 0.535 2.740 0.645 ;
        RECT  2.405 0.535 2.495 1.295 ;
        RECT  2.190 0.535 2.265 0.645 ;
        RECT  2.080 0.535 2.190 1.485 ;
        RECT  2.075 0.535 2.080 0.945 ;
        RECT  2.000 0.775 2.075 0.945 ;
        RECT  1.890 0.535 1.985 0.645 ;
        RECT  1.890 1.045 1.935 1.525 ;
        RECT  1.800 0.535 1.890 1.525 ;
        RECT  0.670 1.435 1.800 1.525 ;
        RECT  1.560 0.275 1.670 1.330 ;
        RECT  1.080 1.235 1.450 1.345 ;
        RECT  1.300 0.340 1.410 0.590 ;
        RECT  1.080 0.500 1.300 0.590 ;
        RECT  0.990 0.500 1.080 1.345 ;
        RECT  0.935 0.500 0.990 0.675 ;
        RECT  0.780 1.235 0.990 1.345 ;
        RECT  0.820 0.265 0.935 0.675 ;
        RECT  0.670 0.780 0.880 0.895 ;
        RECT  0.580 0.575 0.670 1.525 ;
        RECT  0.445 0.575 0.580 0.675 ;
        RECT  0.445 1.425 0.580 1.525 ;
        RECT  0.315 0.265 0.445 0.675 ;
        RECT  0.315 1.040 0.445 1.525 ;
    END
END FCSICIND2

MACRO FCSICOND1
    CLASS CORE ;
    FOREIGN FCSICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.450 0.310 10.550 1.490 ;
        RECT  10.415 0.310 10.450 0.520 ;
        RECT  10.420 1.040 10.450 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0925 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.020 0.700 10.150 1.100 ;
        END
    END CS
    PIN CON1
        ANTENNADIFFAREA 0.1580 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.635 6.165 0.725 ;
        RECT  5.950 1.110 6.150 1.290 ;
        RECT  5.850 0.635 5.950 1.290 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.1580 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.635 5.750 1.290 ;
        RECT  5.445 0.635 5.650 0.725 ;
        RECT  5.450 1.110 5.650 1.290 ;
        END
    END CON0
    PIN CI1
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.640 0.710 8.780 1.090 ;
        END
    END CI1
    PIN CI0
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.710 2.770 1.090 ;
        END
    END CI0
    PIN B
        ANTENNAGATEAREA 0.0927 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.195 0.700 1.350 1.100 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.430 0.895 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 10.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 10.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.330 0.730 10.360 0.940 ;
        RECT  10.240 0.730 10.330 1.525 ;
        RECT  9.455 1.435 10.240 1.525 ;
        RECT  9.930 0.415 10.075 0.525 ;
        RECT  9.930 1.215 10.065 1.345 ;
        RECT  9.830 0.415 9.930 1.345 ;
        RECT  9.750 0.770 9.830 0.940 ;
        RECT  9.660 0.435 9.740 0.625 ;
        RECT  9.660 1.160 9.720 1.345 ;
        RECT  9.570 0.275 9.660 1.345 ;
        RECT  3.590 0.275 9.570 0.365 ;
        RECT  9.455 0.455 9.480 0.625 ;
        RECT  9.345 0.455 9.455 1.525 ;
        RECT  9.080 0.455 9.195 1.495 ;
        RECT  9.055 0.455 9.080 0.665 ;
        RECT  7.875 1.385 9.080 1.495 ;
        RECT  8.475 1.205 8.965 1.295 ;
        RECT  8.475 0.475 8.950 0.565 ;
        RECT  8.365 0.475 8.475 1.295 ;
        RECT  7.750 1.205 8.365 1.295 ;
        RECT  8.090 0.490 8.220 0.600 ;
        RECT  8.000 0.490 8.090 1.115 ;
        RECT  7.875 1.015 8.000 1.115 ;
        RECT  7.800 0.455 7.910 0.875 ;
        RECT  7.750 0.785 7.800 0.875 ;
        RECT  7.650 0.785 7.750 1.295 ;
        RECT  7.560 0.495 7.690 0.605 ;
        RECT  7.470 0.495 7.560 1.295 ;
        RECT  6.615 1.205 7.470 1.295 ;
        RECT  7.270 0.475 7.380 1.115 ;
        RECT  7.055 1.385 7.280 1.500 ;
        RECT  7.065 1.005 7.270 1.115 ;
        RECT  7.075 0.675 7.145 0.885 ;
        RECT  6.975 0.460 7.075 0.885 ;
        RECT  4.555 1.400 7.055 1.500 ;
        RECT  6.965 0.460 6.975 1.115 ;
        RECT  6.885 0.785 6.965 1.115 ;
        RECT  6.805 1.010 6.885 1.115 ;
        RECT  6.705 0.455 6.795 0.900 ;
        RECT  4.905 0.455 6.705 0.545 ;
        RECT  6.525 0.845 6.615 1.295 ;
        RECT  6.455 0.845 6.525 1.015 ;
        RECT  6.365 0.635 6.465 0.725 ;
        RECT  6.365 1.115 6.415 1.295 ;
        RECT  6.275 0.635 6.365 1.295 ;
        RECT  6.060 0.850 6.275 0.980 ;
        RECT  5.335 0.850 5.540 0.980 ;
        RECT  5.245 0.635 5.335 1.295 ;
        RECT  5.125 0.635 5.245 0.725 ;
        RECT  5.195 1.120 5.245 1.295 ;
        RECT  5.085 0.845 5.155 1.015 ;
        RECT  4.995 0.845 5.085 1.295 ;
        RECT  4.150 1.205 4.995 1.295 ;
        RECT  4.815 0.455 4.905 0.900 ;
        RECT  4.725 1.025 4.805 1.115 ;
        RECT  4.650 0.785 4.725 1.115 ;
        RECT  4.635 0.475 4.650 1.115 ;
        RECT  4.475 0.475 4.635 0.895 ;
        RECT  4.330 1.385 4.555 1.500 ;
        RECT  4.350 1.005 4.545 1.115 ;
        RECT  4.240 0.475 4.350 1.115 ;
        RECT  2.190 1.400 4.330 1.500 ;
        RECT  4.060 0.665 4.150 1.295 ;
        RECT  4.040 0.665 4.060 0.755 ;
        RECT  3.930 0.465 4.040 0.755 ;
        RECT  3.860 0.845 3.960 1.295 ;
        RECT  3.790 0.845 3.860 0.935 ;
        RECT  3.050 1.205 3.860 1.295 ;
        RECT  3.680 0.455 3.790 0.935 ;
        RECT  3.590 1.025 3.735 1.115 ;
        RECT  3.500 0.275 3.590 1.115 ;
        RECT  3.380 0.490 3.500 0.600 ;
        RECT  1.670 0.275 3.410 0.380 ;
        RECT  3.290 1.015 3.390 1.115 ;
        RECT  3.200 0.490 3.290 1.115 ;
        RECT  3.105 0.490 3.200 0.600 ;
        RECT  3.015 0.750 3.050 1.295 ;
        RECT  2.925 0.495 3.015 1.295 ;
        RECT  2.550 0.495 2.925 0.605 ;
        RECT  2.550 1.205 2.925 1.295 ;
        RECT  2.190 0.535 2.265 0.645 ;
        RECT  2.080 0.535 2.190 1.500 ;
        RECT  2.075 0.535 2.080 0.945 ;
        RECT  2.000 0.775 2.075 0.945 ;
        RECT  1.890 0.535 1.985 0.645 ;
        RECT  1.890 1.045 1.935 1.525 ;
        RECT  1.800 0.535 1.890 1.525 ;
        RECT  0.670 1.435 1.800 1.525 ;
        RECT  1.560 0.275 1.670 1.330 ;
        RECT  1.080 1.235 1.450 1.345 ;
        RECT  1.300 0.340 1.410 0.590 ;
        RECT  1.080 0.500 1.300 0.590 ;
        RECT  0.990 0.500 1.080 1.345 ;
        RECT  0.935 0.500 0.990 0.675 ;
        RECT  0.780 1.235 0.990 1.345 ;
        RECT  0.820 0.265 0.935 0.675 ;
        RECT  0.670 0.780 0.880 0.895 ;
        RECT  0.580 0.575 0.670 1.525 ;
        RECT  0.445 0.575 0.580 0.675 ;
        RECT  0.445 1.425 0.580 1.525 ;
        RECT  0.315 0.265 0.445 0.675 ;
        RECT  0.315 1.040 0.445 1.525 ;
    END
END FCSICOND1

MACRO FCSICOND2
    CLASS CORE ;
    FOREIGN FCSICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.850 0.275 10.950 1.490 ;
        RECT  10.800 0.275 10.850 0.665 ;
        RECT  10.820 1.040 10.850 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0925 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.420 0.700 10.550 1.100 ;
        END
    END CS
    PIN CON1
        ANTENNADIFFAREA 0.1620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.150 0.635 6.370 0.725 ;
        RECT  6.150 1.110 6.350 1.290 ;
        RECT  6.050 0.635 6.150 1.290 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.1620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.635 5.950 1.290 ;
        RECT  5.640 0.635 5.850 0.725 ;
        RECT  5.650 1.110 5.850 1.290 ;
        END
    END CON0
    PIN CI1
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.040 0.710 9.180 1.090 ;
        END
    END CI1
    PIN CI0
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.710 2.770 1.090 ;
        END
    END CI0
    PIN B
        ANTENNAGATEAREA 0.0927 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.195 0.700 1.350 1.100 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.430 0.895 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 11.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 11.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.730 0.770 10.760 0.940 ;
        RECT  10.640 0.770 10.730 1.525 ;
        RECT  9.855 1.435 10.640 1.525 ;
        RECT  10.330 0.415 10.475 0.525 ;
        RECT  10.330 1.215 10.465 1.345 ;
        RECT  10.230 0.415 10.330 1.345 ;
        RECT  10.150 0.770 10.230 0.940 ;
        RECT  10.060 0.435 10.140 0.625 ;
        RECT  10.060 1.160 10.120 1.345 ;
        RECT  9.970 0.275 10.060 1.345 ;
        RECT  3.590 0.275 9.970 0.365 ;
        RECT  9.855 0.455 9.880 0.625 ;
        RECT  9.745 0.455 9.855 1.525 ;
        RECT  9.480 0.455 9.595 1.495 ;
        RECT  9.455 0.455 9.480 0.665 ;
        RECT  8.275 1.385 9.480 1.495 ;
        RECT  8.875 1.205 9.365 1.295 ;
        RECT  8.875 0.475 9.350 0.565 ;
        RECT  8.765 0.475 8.875 1.295 ;
        RECT  8.150 1.205 8.765 1.295 ;
        RECT  8.490 0.490 8.620 0.600 ;
        RECT  8.400 0.490 8.490 1.115 ;
        RECT  8.275 1.015 8.400 1.115 ;
        RECT  8.200 0.455 8.310 0.875 ;
        RECT  8.150 0.785 8.200 0.875 ;
        RECT  8.050 0.785 8.150 1.295 ;
        RECT  7.960 0.495 8.090 0.605 ;
        RECT  7.870 0.495 7.960 1.295 ;
        RECT  7.015 1.205 7.870 1.295 ;
        RECT  7.670 0.475 7.780 1.115 ;
        RECT  7.455 1.385 7.680 1.500 ;
        RECT  7.465 1.005 7.670 1.115 ;
        RECT  7.475 0.675 7.545 0.885 ;
        RECT  7.375 0.460 7.475 0.885 ;
        RECT  4.535 1.400 7.455 1.500 ;
        RECT  7.365 0.460 7.375 1.115 ;
        RECT  7.285 0.785 7.365 1.115 ;
        RECT  7.205 1.010 7.285 1.115 ;
        RECT  7.105 0.455 7.195 0.900 ;
        RECT  4.905 0.455 7.105 0.545 ;
        RECT  6.925 0.865 7.015 1.295 ;
        RECT  6.775 0.865 6.925 0.995 ;
        RECT  6.665 0.635 6.865 0.735 ;
        RECT  6.665 1.105 6.815 1.295 ;
        RECT  6.555 0.635 6.665 1.295 ;
        RECT  6.240 0.850 6.555 0.980 ;
        RECT  5.455 0.850 5.760 0.980 ;
        RECT  5.345 0.635 5.455 1.295 ;
        RECT  5.125 0.635 5.345 0.735 ;
        RECT  5.195 1.105 5.345 1.295 ;
        RECT  5.085 0.865 5.235 0.995 ;
        RECT  4.995 0.865 5.085 1.295 ;
        RECT  4.150 1.205 4.995 1.295 ;
        RECT  4.815 0.455 4.905 0.900 ;
        RECT  4.725 1.025 4.805 1.115 ;
        RECT  4.650 0.785 4.725 1.115 ;
        RECT  4.635 0.475 4.650 1.115 ;
        RECT  4.475 0.475 4.635 0.895 ;
        RECT  4.350 1.005 4.545 1.115 ;
        RECT  4.325 1.385 4.535 1.500 ;
        RECT  4.240 0.475 4.350 1.115 ;
        RECT  2.190 1.400 4.325 1.500 ;
        RECT  4.060 0.665 4.150 1.295 ;
        RECT  4.040 0.665 4.060 0.755 ;
        RECT  3.930 0.465 4.040 0.755 ;
        RECT  3.860 0.845 3.960 1.295 ;
        RECT  3.790 0.845 3.860 0.935 ;
        RECT  3.050 1.205 3.860 1.295 ;
        RECT  3.680 0.455 3.790 0.935 ;
        RECT  3.590 1.025 3.735 1.115 ;
        RECT  3.500 0.275 3.590 1.115 ;
        RECT  3.380 0.490 3.500 0.600 ;
        RECT  1.670 0.275 3.410 0.380 ;
        RECT  3.290 1.015 3.390 1.115 ;
        RECT  3.200 0.490 3.290 1.115 ;
        RECT  3.105 0.490 3.200 0.600 ;
        RECT  3.015 0.750 3.050 1.295 ;
        RECT  2.925 0.495 3.015 1.295 ;
        RECT  2.550 0.495 2.925 0.605 ;
        RECT  2.550 1.205 2.925 1.295 ;
        RECT  2.190 0.535 2.265 0.645 ;
        RECT  2.080 0.535 2.190 1.500 ;
        RECT  2.075 0.535 2.080 0.945 ;
        RECT  2.000 0.775 2.075 0.945 ;
        RECT  1.890 0.535 1.985 0.645 ;
        RECT  1.890 1.045 1.935 1.525 ;
        RECT  1.800 0.535 1.890 1.525 ;
        RECT  0.670 1.435 1.800 1.525 ;
        RECT  1.560 0.275 1.670 1.330 ;
        RECT  1.080 1.235 1.450 1.345 ;
        RECT  1.300 0.340 1.410 0.590 ;
        RECT  1.080 0.500 1.300 0.590 ;
        RECT  0.990 0.500 1.080 1.345 ;
        RECT  0.935 0.500 0.990 0.675 ;
        RECT  0.780 1.235 0.990 1.345 ;
        RECT  0.820 0.265 0.935 0.675 ;
        RECT  0.670 0.780 0.880 0.895 ;
        RECT  0.580 0.575 0.670 1.525 ;
        RECT  0.445 0.575 0.580 0.675 ;
        RECT  0.445 1.425 0.580 1.525 ;
        RECT  0.315 0.265 0.445 0.675 ;
        RECT  0.315 1.040 0.445 1.525 ;
    END
END FCSICOND2

MACRO FICIND1
    CLASS CORE ;
    FOREIGN FICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.625 0.275 5.750 1.490 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.150 0.425 5.245 0.535 ;
        RECT  5.150 1.015 5.245 1.115 ;
        RECT  5.050 0.425 5.150 1.115 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0527 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.710 4.390 0.890 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.0927 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.550 0.890 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.460 -0.165 5.800 0.165 ;
        RECT  5.350 -0.165 5.460 0.585 ;
        RECT  1.305 -0.165 5.350 0.165 ;
        RECT  1.135 -0.165 1.305 0.410 ;
        RECT  0.785 -0.165 1.135 0.165 ;
        RECT  0.615 -0.165 0.785 0.420 ;
        RECT  0.235 -0.165 0.615 0.165 ;
        RECT  0.125 -0.165 0.235 0.585 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.510 1.635 5.800 1.965 ;
        RECT  5.400 1.385 5.510 1.965 ;
        RECT  5.300 1.385 5.400 1.495 ;
        RECT  1.330 1.635 5.400 1.965 ;
        RECT  1.140 1.505 1.330 1.965 ;
        RECT  0.705 1.635 1.140 1.965 ;
        RECT  0.705 1.385 0.805 1.495 ;
        RECT  0.595 1.385 0.705 1.965 ;
        RECT  0.235 1.635 0.595 1.965 ;
        RECT  0.125 1.040 0.235 1.965 ;
        RECT  0.000 1.635 0.125 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.430 0.730 5.535 1.295 ;
        RECT  3.960 1.205 5.430 1.295 ;
        RECT  3.395 1.430 5.080 1.520 ;
        RECT  4.850 0.475 4.940 1.115 ;
        RECT  4.810 0.475 4.850 0.585 ;
        RECT  4.715 1.015 4.850 1.115 ;
        RECT  4.715 0.275 4.810 0.585 ;
        RECT  4.600 0.755 4.740 0.865 ;
        RECT  3.770 0.275 4.715 0.365 ;
        RECT  4.590 0.755 4.600 1.115 ;
        RECT  4.500 0.455 4.590 1.115 ;
        RECT  4.160 0.455 4.500 0.565 ;
        RECT  4.050 1.005 4.500 1.115 ;
        RECT  3.960 0.500 4.070 0.610 ;
        RECT  3.870 0.500 3.960 1.295 ;
        RECT  3.755 1.185 3.870 1.295 ;
        RECT  3.660 0.275 3.770 0.880 ;
        RECT  3.655 0.790 3.660 0.880 ;
        RECT  3.545 0.790 3.655 1.330 ;
        RECT  3.395 0.485 3.535 0.595 ;
        RECT  3.280 0.485 3.395 1.520 ;
        RECT  3.100 0.435 3.190 1.470 ;
        RECT  2.350 1.360 3.100 1.470 ;
        RECT  2.900 0.595 3.010 1.250 ;
        RECT  2.895 0.595 2.900 0.695 ;
        RECT  2.710 1.140 2.900 1.250 ;
        RECT  2.785 0.275 2.895 0.695 ;
        RECT  2.640 0.785 2.780 0.890 ;
        RECT  2.550 0.285 2.640 0.890 ;
        RECT  1.830 0.285 2.550 0.375 ;
        RECT  2.350 0.465 2.425 0.575 ;
        RECT  2.235 0.465 2.350 1.470 ;
        RECT  2.160 0.775 2.235 0.945 ;
        RECT  2.050 0.465 2.145 0.575 ;
        RECT  2.050 1.060 2.095 1.525 ;
        RECT  1.960 0.465 2.050 1.525 ;
        RECT  1.530 1.435 1.960 1.525 ;
        RECT  1.720 0.285 1.830 1.325 ;
        RECT  1.160 0.500 1.620 0.600 ;
        RECT  1.320 1.125 1.620 1.235 ;
        RECT  1.440 1.325 1.530 1.525 ;
        RECT  1.045 1.325 1.440 1.415 ;
        RECT  1.230 1.015 1.320 1.235 ;
        RECT  1.160 1.015 1.230 1.115 ;
        RECT  1.070 0.500 1.160 1.115 ;
        RECT  1.015 0.500 1.070 0.695 ;
        RECT  0.855 1.005 1.070 1.115 ;
        RECT  0.955 1.205 1.045 1.415 ;
        RECT  0.900 0.275 1.015 0.695 ;
        RECT  0.750 0.785 0.960 0.895 ;
        RECT  0.750 1.205 0.955 1.295 ;
        RECT  0.660 0.530 0.750 1.295 ;
        RECT  0.495 0.530 0.660 0.620 ;
        RECT  0.495 1.205 0.660 1.295 ;
        RECT  0.385 0.375 0.495 0.620 ;
        RECT  0.385 1.040 0.495 1.470 ;
    END
END FICIND1

MACRO FICIND2
    CLASS CORE ;
    FOREIGN FICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.310 5.950 1.325 ;
        RECT  5.835 0.310 5.850 0.585 ;
        RECT  5.835 1.115 5.850 1.325 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.475 0.570 6.550 1.150 ;
        RECT  6.450 0.275 6.475 1.470 ;
        RECT  6.345 0.275 6.450 0.695 ;
        RECT  6.345 1.040 6.450 1.470 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.710 4.950 0.890 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.1483 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.645 0.710 2.755 1.090 ;
        RECT  2.610 0.710 2.645 0.895 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 -0.165 6.800 0.165 ;
        RECT  6.615 -0.165 6.725 0.455 ;
        RECT  6.205 -0.165 6.615 0.165 ;
        RECT  6.095 -0.165 6.205 0.695 ;
        RECT  5.685 -0.165 6.095 0.165 ;
        RECT  5.575 -0.165 5.685 0.585 ;
        RECT  0.785 -0.165 5.575 0.165 ;
        RECT  0.615 -0.165 0.785 0.420 ;
        RECT  0.235 -0.165 0.615 0.165 ;
        RECT  0.125 -0.165 0.235 0.585 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 1.635 6.800 1.965 ;
        RECT  6.615 1.260 6.725 1.965 ;
        RECT  0.785 1.635 6.615 1.965 ;
        RECT  0.615 1.385 0.785 1.965 ;
        RECT  0.235 1.635 0.615 1.965 ;
        RECT  0.125 1.040 0.235 1.965 ;
        RECT  0.000 1.635 0.125 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.215 0.785 6.340 0.895 ;
        RECT  6.105 0.785 6.215 1.525 ;
        RECT  3.555 1.435 6.105 1.525 ;
        RECT  5.685 0.750 5.760 0.920 ;
        RECT  5.575 0.750 5.685 1.345 ;
        RECT  4.105 1.255 5.575 1.345 ;
        RECT  5.335 0.275 5.430 1.165 ;
        RECT  5.320 0.275 5.335 0.655 ;
        RECT  5.320 0.995 5.335 1.165 ;
        RECT  3.920 0.275 5.320 0.365 ;
        RECT  5.180 0.740 5.245 0.910 ;
        RECT  5.070 0.480 5.180 1.165 ;
        RECT  4.285 0.480 5.070 0.615 ;
        RECT  4.215 1.055 5.070 1.165 ;
        RECT  4.105 0.455 4.175 0.890 ;
        RECT  4.060 0.455 4.105 1.345 ;
        RECT  4.015 0.780 4.060 1.345 ;
        RECT  3.925 1.185 4.015 1.345 ;
        RECT  3.815 0.275 3.920 1.035 ;
        RECT  3.805 0.275 3.815 1.290 ;
        RECT  3.695 0.945 3.805 1.290 ;
        RECT  3.555 0.445 3.645 0.840 ;
        RECT  3.535 0.445 3.555 1.525 ;
        RECT  3.445 0.725 3.535 1.525 ;
        RECT  3.350 0.505 3.415 0.615 ;
        RECT  3.245 0.505 3.350 1.470 ;
        RECT  2.035 0.275 3.295 0.385 ;
        RECT  2.555 1.355 3.245 1.470 ;
        RECT  3.045 0.535 3.155 1.135 ;
        RECT  2.920 0.535 3.045 0.645 ;
        RECT  2.920 1.025 3.045 1.135 ;
        RECT  2.520 0.495 2.630 0.595 ;
        RECT  2.520 1.005 2.555 1.470 ;
        RECT  2.420 0.495 2.520 1.470 ;
        RECT  2.325 0.775 2.420 0.945 ;
        RECT  2.235 0.475 2.310 0.645 ;
        RECT  2.235 1.060 2.295 1.525 ;
        RECT  2.145 0.475 2.235 1.525 ;
        RECT  1.005 1.435 2.145 1.525 ;
        RECT  1.925 0.275 2.035 1.325 ;
        RECT  1.245 1.235 1.825 1.345 ;
        RECT  1.665 0.275 1.775 0.535 ;
        RECT  1.545 0.780 1.670 0.890 ;
        RECT  1.245 0.275 1.665 0.365 ;
        RECT  1.525 0.780 1.545 1.125 ;
        RECT  1.355 0.475 1.525 1.125 ;
        RECT  1.155 0.275 1.245 1.345 ;
        RECT  1.015 0.585 1.155 0.695 ;
        RECT  0.855 1.005 1.155 1.115 ;
        RECT  0.750 0.785 1.045 0.895 ;
        RECT  0.900 0.275 1.015 0.695 ;
        RECT  0.915 1.205 1.005 1.525 ;
        RECT  0.750 1.205 0.915 1.295 ;
        RECT  0.660 0.530 0.750 1.295 ;
        RECT  0.495 0.530 0.660 0.620 ;
        RECT  0.495 1.205 0.660 1.295 ;
        RECT  0.385 0.375 0.495 0.620 ;
        RECT  0.385 1.040 0.495 1.470 ;
    END
END FICIND2

MACRO FICOND1
    CLASS CORE ;
    FOREIGN FICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.025 0.275 6.150 1.490 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.1400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.510 5.750 1.115 ;
        RECT  5.540 0.275 5.650 0.695 ;
        RECT  5.500 1.005 5.650 1.115 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0445 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.710 4.950 0.890 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0927 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.550 0.890 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 -0.165 6.200 0.165 ;
        RECT  1.135 -0.165 1.305 0.410 ;
        RECT  0.785 -0.165 1.135 0.165 ;
        RECT  0.615 -0.165 0.785 0.420 ;
        RECT  0.235 -0.165 0.615 0.165 ;
        RECT  0.125 -0.165 0.235 0.585 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.635 6.200 1.965 ;
        RECT  1.140 1.505 1.330 1.965 ;
        RECT  0.785 1.635 1.140 1.965 ;
        RECT  0.615 1.385 0.785 1.965 ;
        RECT  0.235 1.635 0.615 1.965 ;
        RECT  0.125 1.040 0.235 1.965 ;
        RECT  0.000 1.635 0.125 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.840 0.730 5.935 1.295 ;
        RECT  3.960 1.205 5.840 1.295 ;
        RECT  5.310 0.785 5.555 0.895 ;
        RECT  5.200 0.585 5.310 1.115 ;
        RECT  5.150 0.585 5.200 0.695 ;
        RECT  5.000 1.005 5.200 1.115 ;
        RECT  5.040 0.275 5.150 0.695 ;
        RECT  3.395 1.430 5.045 1.520 ;
        RECT  4.515 0.475 4.910 0.585 ;
        RECT  4.515 1.005 4.910 1.115 ;
        RECT  4.405 0.275 4.515 1.115 ;
        RECT  3.770 0.275 4.405 0.365 ;
        RECT  4.190 0.455 4.300 1.115 ;
        RECT  4.050 1.005 4.190 1.115 ;
        RECT  3.960 0.500 4.070 0.610 ;
        RECT  3.870 0.500 3.960 1.295 ;
        RECT  3.755 1.185 3.870 1.295 ;
        RECT  3.660 0.275 3.770 0.880 ;
        RECT  3.655 0.790 3.660 0.880 ;
        RECT  3.545 0.790 3.655 1.330 ;
        RECT  3.395 0.485 3.535 0.595 ;
        RECT  3.280 0.485 3.395 1.520 ;
        RECT  3.100 0.435 3.190 1.470 ;
        RECT  2.350 1.360 3.100 1.470 ;
        RECT  2.900 0.595 3.010 1.250 ;
        RECT  2.895 0.595 2.900 0.695 ;
        RECT  2.710 1.140 2.900 1.250 ;
        RECT  2.785 0.275 2.895 0.695 ;
        RECT  2.640 0.785 2.780 0.890 ;
        RECT  2.550 0.285 2.640 0.890 ;
        RECT  1.830 0.285 2.550 0.375 ;
        RECT  2.350 0.465 2.425 0.575 ;
        RECT  2.235 0.465 2.350 1.470 ;
        RECT  2.160 0.775 2.235 0.945 ;
        RECT  2.050 0.465 2.145 0.575 ;
        RECT  2.050 1.060 2.095 1.525 ;
        RECT  1.960 0.465 2.050 1.525 ;
        RECT  1.530 1.435 1.960 1.525 ;
        RECT  1.720 0.285 1.830 1.325 ;
        RECT  1.160 0.500 1.620 0.600 ;
        RECT  1.320 1.125 1.620 1.235 ;
        RECT  1.440 1.325 1.530 1.525 ;
        RECT  1.045 1.325 1.440 1.415 ;
        RECT  1.230 1.015 1.320 1.235 ;
        RECT  1.160 1.015 1.230 1.115 ;
        RECT  1.070 0.500 1.160 1.115 ;
        RECT  1.015 0.500 1.070 0.695 ;
        RECT  0.855 1.005 1.070 1.115 ;
        RECT  0.955 1.205 1.045 1.415 ;
        RECT  0.900 0.275 1.015 0.695 ;
        RECT  0.750 0.785 0.960 0.895 ;
        RECT  0.750 1.205 0.955 1.295 ;
        RECT  0.660 0.530 0.750 1.295 ;
        RECT  0.495 0.530 0.660 0.620 ;
        RECT  0.495 1.205 0.660 1.295 ;
        RECT  0.385 0.375 0.495 0.620 ;
        RECT  0.385 1.040 0.495 1.470 ;
    END
END FICOND1

MACRO FICOND2
    CLASS CORE ;
    FOREIGN FICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.475 0.570 6.550 1.150 ;
        RECT  6.450 0.275 6.475 1.470 ;
        RECT  6.345 0.275 6.450 0.695 ;
        RECT  6.345 1.040 6.450 1.470 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.845 0.275 5.950 1.165 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 5.160 0.890 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.1483 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.645 0.710 2.755 1.090 ;
        RECT  2.610 0.710 2.645 0.895 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 -0.165 6.800 0.165 ;
        RECT  6.615 -0.165 6.725 0.455 ;
        RECT  6.205 -0.165 6.615 0.165 ;
        RECT  6.095 -0.165 6.205 0.695 ;
        RECT  5.685 -0.165 6.095 0.165 ;
        RECT  5.575 -0.165 5.685 0.585 ;
        RECT  0.785 -0.165 5.575 0.165 ;
        RECT  0.615 -0.165 0.785 0.420 ;
        RECT  0.235 -0.165 0.615 0.165 ;
        RECT  0.125 -0.165 0.235 0.585 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 1.635 6.800 1.965 ;
        RECT  6.615 1.260 6.725 1.965 ;
        RECT  0.785 1.635 6.615 1.965 ;
        RECT  0.615 1.385 0.785 1.965 ;
        RECT  0.235 1.635 0.615 1.965 ;
        RECT  0.125 1.040 0.235 1.965 ;
        RECT  0.000 1.635 0.125 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.215 0.785 6.340 0.895 ;
        RECT  6.105 0.785 6.215 1.345 ;
        RECT  4.105 1.255 6.105 1.345 ;
        RECT  5.425 0.750 5.755 0.920 ;
        RECT  5.330 1.435 5.540 1.545 ;
        RECT  5.295 0.275 5.425 1.165 ;
        RECT  3.555 1.435 5.330 1.525 ;
        RECT  4.605 0.400 4.985 0.535 ;
        RECT  4.605 1.055 4.985 1.165 ;
        RECT  4.515 0.275 4.605 1.165 ;
        RECT  3.920 0.275 4.515 0.365 ;
        RECT  4.490 0.730 4.515 0.900 ;
        RECT  4.400 0.455 4.425 0.625 ;
        RECT  4.285 0.455 4.400 1.165 ;
        RECT  4.215 1.055 4.285 1.165 ;
        RECT  4.105 0.455 4.175 0.890 ;
        RECT  4.060 0.455 4.105 1.345 ;
        RECT  4.015 0.780 4.060 1.345 ;
        RECT  3.925 1.185 4.015 1.345 ;
        RECT  3.815 0.275 3.920 1.035 ;
        RECT  3.805 0.275 3.815 1.290 ;
        RECT  3.695 0.945 3.805 1.290 ;
        RECT  3.555 0.445 3.645 0.840 ;
        RECT  3.535 0.445 3.555 1.525 ;
        RECT  3.445 0.725 3.535 1.525 ;
        RECT  3.350 0.505 3.415 0.615 ;
        RECT  3.245 0.505 3.350 1.470 ;
        RECT  2.035 0.275 3.295 0.385 ;
        RECT  2.555 1.355 3.245 1.470 ;
        RECT  3.045 0.535 3.155 1.135 ;
        RECT  2.920 0.535 3.045 0.645 ;
        RECT  2.920 1.025 3.045 1.135 ;
        RECT  2.520 0.495 2.630 0.595 ;
        RECT  2.520 1.005 2.555 1.470 ;
        RECT  2.420 0.495 2.520 1.470 ;
        RECT  2.325 0.775 2.420 0.945 ;
        RECT  2.235 0.475 2.310 0.645 ;
        RECT  2.235 1.060 2.295 1.525 ;
        RECT  2.145 0.475 2.235 1.525 ;
        RECT  1.005 1.435 2.145 1.525 ;
        RECT  1.925 0.275 2.035 1.325 ;
        RECT  1.245 1.235 1.825 1.345 ;
        RECT  1.665 0.275 1.775 0.535 ;
        RECT  1.545 0.780 1.670 0.890 ;
        RECT  1.245 0.275 1.665 0.365 ;
        RECT  1.525 0.780 1.545 1.125 ;
        RECT  1.355 0.475 1.525 1.125 ;
        RECT  1.155 0.275 1.245 1.345 ;
        RECT  1.015 0.585 1.155 0.695 ;
        RECT  0.855 1.005 1.155 1.115 ;
        RECT  0.750 0.785 1.045 0.895 ;
        RECT  0.900 0.275 1.015 0.695 ;
        RECT  0.915 1.205 1.005 1.525 ;
        RECT  0.750 1.205 0.915 1.295 ;
        RECT  0.660 0.530 0.750 1.295 ;
        RECT  0.495 0.530 0.660 0.620 ;
        RECT  0.495 1.205 0.660 1.295 ;
        RECT  0.385 0.375 0.495 0.620 ;
        RECT  0.385 1.040 0.495 1.470 ;
    END
END FICOND2

MACRO FIICOND1
    CLASS CORE ;
    FOREIGN FIICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.275 5.750 1.490 ;
        RECT  5.615 0.275 5.650 0.665 ;
        RECT  5.615 1.040 5.650 1.490 ;
        END
    END S
    PIN CON1
        ANTENNADIFFAREA 0.1530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.090 1.195 1.200 ;
        RECT  0.850 0.490 0.970 1.200 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.1660 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 1.200 0.455 1.455 ;
        RECT  0.150 1.200 0.315 1.290 ;
        RECT  0.150 0.310 0.175 0.520 ;
        RECT  0.050 0.310 0.150 1.290 ;
        END
    END CON0
    PIN C
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.045 0.700 5.155 1.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.2029 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.425 3.255 1.525 ;
        RECT  1.050 1.375 1.150 1.525 ;
        RECT  0.750 1.375 1.050 1.465 ;
        RECT  0.650 0.710 0.750 1.465 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.2204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.780 1.550 0.890 ;
        RECT  1.110 0.290 1.210 0.890 ;
        RECT  0.375 0.290 1.110 0.380 ;
        RECT  0.265 0.290 0.375 1.090 ;
        RECT  0.250 0.705 0.265 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.465 1.635 5.800 1.965 ;
        RECT  5.355 1.055 5.465 1.965 ;
        RECT  0.000 1.635 5.355 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.525 0.755 5.560 0.945 ;
        RECT  5.425 0.275 5.525 0.945 ;
        RECT  4.440 0.275 5.425 0.365 ;
        RECT  4.905 0.480 5.275 0.590 ;
        RECT  4.905 1.210 5.255 1.320 ;
        RECT  4.815 0.480 4.905 1.525 ;
        RECT  4.755 0.755 4.815 0.925 ;
        RECT  4.155 1.435 4.815 1.525 ;
        RECT  4.665 0.455 4.725 0.645 ;
        RECT  4.565 0.455 4.665 1.345 ;
        RECT  4.415 0.275 4.440 0.645 ;
        RECT  4.330 0.275 4.415 1.345 ;
        RECT  4.305 0.515 4.330 1.345 ;
        RECT  3.920 0.285 4.220 0.415 ;
        RECT  4.045 0.515 4.155 1.525 ;
        RECT  3.820 0.285 3.920 1.470 ;
        RECT  3.785 0.285 3.820 0.665 ;
        RECT  3.785 1.040 3.820 1.470 ;
        RECT  3.645 0.750 3.730 0.920 ;
        RECT  3.555 0.750 3.645 1.335 ;
        RECT  2.860 1.245 3.555 1.335 ;
        RECT  3.285 0.275 3.395 1.155 ;
        RECT  3.165 0.750 3.285 0.920 ;
        RECT  3.050 0.310 3.175 0.420 ;
        RECT  3.050 1.025 3.170 1.135 ;
        RECT  2.960 0.310 3.050 1.135 ;
        RECT  1.795 0.310 2.960 0.400 ;
        RECT  2.835 0.810 2.860 1.335 ;
        RECT  2.750 0.510 2.835 1.335 ;
        RECT  2.725 0.510 2.750 0.900 ;
        RECT  2.490 0.510 2.605 1.325 ;
        RECT  1.905 0.510 2.490 0.620 ;
        RECT  1.965 1.215 2.490 1.325 ;
        RECT  1.795 0.780 2.145 0.890 ;
        RECT  1.700 0.310 1.795 1.325 ;
        RECT  1.520 0.565 1.700 0.665 ;
        RECT  1.465 1.215 1.700 1.325 ;
        RECT  1.410 0.275 1.520 0.665 ;
    END
END FIICOND1

MACRO FIICOND2
    CLASS CORE ;
    FOREIGN FIICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.565 6.750 1.140 ;
        RECT  6.540 0.275 6.650 0.665 ;
        RECT  6.540 1.040 6.650 1.470 ;
        END
    END S
    PIN CON1
        ANTENNADIFFAREA 0.2600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.860 0.510 2.015 0.620 ;
        RECT  1.770 0.510 1.860 1.300 ;
        RECT  1.465 1.100 1.770 1.300 ;
        RECT  1.355 0.490 1.465 1.300 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.2860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.205 0.985 1.315 ;
        RECT  0.585 0.275 0.750 0.675 ;
        RECT  0.550 0.575 0.585 0.675 ;
        RECT  0.450 0.575 0.550 1.315 ;
        RECT  0.250 1.205 0.450 1.315 ;
        END
    END CON0
    PIN C
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.045 0.700 6.155 1.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.3130 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.425 4.180 1.525 ;
        RECT  1.950 0.730 2.050 1.525 ;
        RECT  1.200 1.425 1.950 1.525 ;
        RECT  1.090 0.710 1.200 1.525 ;
        RECT  0.150 1.425 1.090 1.525 ;
        RECT  0.150 0.780 0.350 0.890 ;
        RECT  0.050 0.780 0.150 1.525 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.3302 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.780 2.475 0.890 ;
        RECT  2.145 0.290 2.245 0.890 ;
        RECT  1.680 0.290 2.145 0.380 ;
        RECT  1.570 0.290 1.680 0.930 ;
        RECT  0.970 0.290 1.570 0.380 ;
        RECT  0.850 0.290 0.970 0.890 ;
        RECT  0.690 0.775 0.850 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.910 -0.165 7.000 0.165 ;
        RECT  6.800 -0.165 6.910 0.465 ;
        RECT  0.195 -0.165 6.800 0.165 ;
        RECT  0.085 -0.165 0.195 0.690 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.910 1.635 7.000 1.965 ;
        RECT  6.800 1.355 6.910 1.965 ;
        RECT  6.390 1.635 6.800 1.965 ;
        RECT  6.280 1.055 6.390 1.965 ;
        RECT  0.000 1.635 6.280 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.430 0.785 6.550 0.895 ;
        RECT  6.330 0.275 6.430 0.895 ;
        RECT  5.365 0.275 6.330 0.365 ;
        RECT  5.830 0.480 6.200 0.590 ;
        RECT  5.830 1.210 6.180 1.320 ;
        RECT  5.740 0.480 5.830 1.525 ;
        RECT  5.680 0.755 5.740 0.925 ;
        RECT  5.080 1.435 5.740 1.525 ;
        RECT  5.590 0.455 5.650 0.645 ;
        RECT  5.490 0.455 5.590 1.345 ;
        RECT  5.340 0.275 5.365 0.645 ;
        RECT  5.255 0.275 5.340 1.345 ;
        RECT  5.230 0.515 5.255 1.345 ;
        RECT  5.080 0.465 5.125 1.140 ;
        RECT  5.015 0.465 5.080 1.525 ;
        RECT  4.970 0.465 5.015 0.655 ;
        RECT  4.970 1.030 5.015 1.525 ;
        RECT  4.845 0.750 4.925 0.920 ;
        RECT  4.745 0.285 4.845 1.470 ;
        RECT  4.710 0.285 4.745 0.665 ;
        RECT  4.710 1.040 4.745 1.470 ;
        RECT  4.570 0.750 4.655 0.920 ;
        RECT  4.480 0.750 4.570 1.335 ;
        RECT  3.785 1.245 4.480 1.335 ;
        RECT  4.210 0.275 4.320 1.155 ;
        RECT  4.090 0.750 4.210 0.920 ;
        RECT  3.975 0.310 4.100 0.420 ;
        RECT  3.975 1.025 4.095 1.135 ;
        RECT  3.885 0.310 3.975 1.135 ;
        RECT  2.720 0.310 3.885 0.400 ;
        RECT  3.760 0.810 3.785 1.335 ;
        RECT  3.675 0.510 3.760 1.335 ;
        RECT  3.650 0.510 3.675 0.900 ;
        RECT  3.415 0.510 3.530 1.325 ;
        RECT  2.830 0.510 3.415 0.620 ;
        RECT  2.850 1.215 3.415 1.325 ;
        RECT  2.720 0.780 3.070 0.890 ;
        RECT  2.625 0.310 2.720 1.325 ;
        RECT  2.465 0.565 2.625 0.665 ;
        RECT  2.310 1.215 2.625 1.325 ;
        RECT  2.355 0.275 2.465 0.665 ;
    END
END FIICOND2

MACRO FILL1
    CLASS CORE ;
    FOREIGN FILL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 0.200 1.965 ;
        END
    END VDD
END FILL1

MACRO FILL16
    CLASS CORE ;
    FOREIGN FILL16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.200 1.965 ;
        END
    END VDD
END FILL16

MACRO FILL1_LL
    CLASS CORE ;
    FOREIGN FILL1_LL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 0.200 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.000 0.310 0.200 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.200 0.165 ;
        RECT  0.000 3.435 0.200 3.765 ;
        END
    END VDD
END FILL1_LL

MACRO FILL2
    CLASS CORE ;
    FOREIGN FILL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 0.400 1.965 ;
        END
    END VDD
END FILL2

MACRO FILL32
    CLASS CORE ;
    FOREIGN FILL32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 6.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 6.400 1.965 ;
        END
    END VDD
END FILL32

MACRO FILL4
    CLASS CORE ;
    FOREIGN FILL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 0.800 1.965 ;
        END
    END VDD
END FILL4

MACRO FILL64
    CLASS CORE ;
    FOREIGN FILL64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 12.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 12.800 1.965 ;
        END
    END VDD
END FILL64

MACRO FILL8
    CLASS CORE ;
    FOREIGN FILL8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VDD
END FILL8

MACRO FILL_NW_HH
    CLASS CORE ;
    FOREIGN FILL_NW_HH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        RECT  0.000 3.435 1.600 3.765 ;
        END
    END VDD
END FILL_NW_HH

MACRO FILL_NW_LL
    CLASS CORE ;
    FOREIGN FILL_NW_LL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.200 -0.165 1.600 0.165 ;
        RECT  1.200 3.435 1.600 3.765 ;
        END
    END VDD
END FILL_NW_LL

MACRO GAN2D1
    CLASS CORE ;
    FOREIGN GAN2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 0.495 1.550 1.525 ;
        RECT  1.450 0.275 1.515 1.525 ;
        RECT  1.405 0.275 1.450 0.585 ;
        RECT  1.405 1.240 1.450 1.525 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.690 0.350 1.095 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.095 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.025 -0.165 1.600 0.165 ;
        RECT  1.025 0.305 1.285 0.415 ;
        RECT  0.855 -0.165 1.025 0.415 ;
        RECT  0.195 -0.165 0.855 0.165 ;
        RECT  0.085 -0.165 0.195 0.455 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.995 1.635 1.600 1.965 ;
        RECT  0.995 1.210 1.285 1.320 ;
        RECT  0.885 1.210 0.995 1.965 ;
        RECT  0.745 1.635 0.885 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.195 1.635 0.575 1.965 ;
        RECT  0.085 1.335 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.730 1.360 1.110 ;
        RECT  0.760 1.000 1.250 1.110 ;
        RECT  0.940 0.610 1.140 0.910 ;
        RECT  0.715 0.470 0.760 1.305 ;
        RECT  0.660 0.275 0.715 1.305 ;
        RECT  0.605 0.275 0.660 0.580 ;
        RECT  0.315 1.205 0.660 1.305 ;
        RECT  0.315 0.275 0.485 0.580 ;
    END
END GAN2D1

MACRO GAN2D2
    CLASS CORE ;
    FOREIGN GAN2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.305 ;
        RECT  1.255 0.510 1.450 0.610 ;
        RECT  1.115 1.205 1.450 1.305 ;
        RECT  1.145 0.275 1.255 0.610 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.690 0.350 1.095 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.095 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  0.995 -0.165 1.375 0.165 ;
        RECT  0.885 -0.165 0.995 0.465 ;
        RECT  0.195 -0.165 0.885 0.165 ;
        RECT  0.085 -0.165 0.195 0.455 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.635 1.600 1.965 ;
        RECT  1.375 1.395 1.545 1.965 ;
        RECT  0.995 1.635 1.375 1.965 ;
        RECT  0.885 1.335 0.995 1.965 ;
        RECT  0.745 1.635 0.885 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.195 1.635 0.575 1.965 ;
        RECT  0.085 1.335 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.730 1.360 1.110 ;
        RECT  1.140 1.000 1.250 1.110 ;
        RECT  1.030 0.730 1.140 1.110 ;
        RECT  0.760 1.000 1.030 1.110 ;
        RECT  0.715 0.470 0.760 1.305 ;
        RECT  0.660 0.275 0.715 1.305 ;
        RECT  0.605 0.275 0.660 0.580 ;
        RECT  0.315 1.205 0.660 1.305 ;
        RECT  0.315 0.275 0.485 0.580 ;
    END
END GAN2D2

MACRO GAOI21D1
    CLASS CORE ;
    FOREIGN GAOI21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.275 1.005 0.490 ;
        RECT  0.650 0.275 0.750 1.305 ;
        RECT  0.595 0.275 0.650 0.445 ;
        RECT  0.315 1.205 0.650 1.305 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.690 1.150 1.095 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.690 0.350 1.095 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.095 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.415 ;
        RECT  0.195 -0.165 1.375 0.165 ;
        RECT  1.115 0.305 1.375 0.415 ;
        RECT  0.085 -0.165 0.195 0.455 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.210 1.515 1.965 ;
        RECT  1.115 1.210 1.405 1.320 ;
        RECT  0.000 1.635 1.405 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.610 1.460 0.910 ;
        RECT  0.885 1.335 0.995 1.525 ;
        RECT  0.195 1.395 0.885 1.525 ;
        RECT  0.315 0.275 0.485 0.580 ;
        RECT  0.085 1.335 0.195 1.525 ;
    END
END GAOI21D1

MACRO GAOI21D2
    CLASS CORE ;
    FOREIGN GAOI21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.4720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.315 0.495 2.350 1.305 ;
        RECT  2.250 0.275 2.315 1.305 ;
        RECT  2.205 0.275 2.250 0.600 ;
        RECT  0.950 1.205 2.250 1.305 ;
        RECT  0.950 0.275 0.995 0.585 ;
        RECT  0.885 0.275 0.950 1.305 ;
        RECT  0.850 0.495 0.885 1.305 ;
        RECT  0.715 0.495 0.850 0.585 ;
        RECT  0.605 0.275 0.715 0.585 ;
        RECT  0.195 0.495 0.605 0.585 ;
        RECT  0.050 0.275 0.195 0.585 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.695 0.560 1.095 ;
        RECT  0.350 0.985 0.450 1.095 ;
        RECT  0.240 0.695 0.350 1.095 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.695 1.950 0.910 ;
        RECT  1.360 0.800 1.840 0.910 ;
        RECT  1.250 0.695 1.360 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.695 2.160 1.115 ;
        RECT  1.150 1.020 2.050 1.115 ;
        RECT  1.040 0.695 1.150 1.115 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.825 -0.165 2.400 0.165 ;
        RECT  1.655 -0.165 1.825 0.405 ;
        RECT  1.545 -0.165 1.655 0.165 ;
        RECT  1.375 -0.165 1.545 0.405 ;
        RECT  0.485 -0.165 1.375 0.165 ;
        RECT  0.315 -0.165 0.485 0.405 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 1.635 2.400 1.965 ;
        RECT  0.315 1.205 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 1.395 2.345 1.525 ;
        RECT  1.935 0.275 2.095 0.585 ;
        RECT  1.105 0.275 1.265 0.585 ;
        RECT  0.575 1.210 0.750 1.525 ;
        RECT  0.050 1.210 0.225 1.525 ;
        LAYER VIA1 ;
        RECT  0.650 1.350 0.750 1.450 ;
        RECT  0.090 1.350 0.190 1.450 ;
        LAYER M2 ;
        RECT  0.650 1.310 0.750 1.490 ;
        RECT  0.150 1.350 0.650 1.450 ;
        RECT  0.050 1.310 0.150 1.490 ;
    END
END GAOI21D2

MACRO GAOI22D1
    CLASS CORE ;
    FOREIGN GAOI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.560 1.550 1.500 ;
        RECT  1.340 0.560 1.450 0.650 ;
        RECT  0.845 1.390 1.450 1.500 ;
        RECT  1.240 0.530 1.340 0.650 ;
        RECT  0.985 0.530 1.240 0.620 ;
        RECT  0.875 0.275 0.985 0.620 ;
        RECT  0.850 0.275 0.875 0.530 ;
        RECT  0.750 0.440 0.850 0.530 ;
        RECT  0.605 0.275 0.750 0.530 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.690 0.350 1.095 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.095 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.740 1.360 1.100 ;
        RECT  0.750 1.010 1.250 1.100 ;
        RECT  0.650 0.690 0.750 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 1.150 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.165 1.600 0.165 ;
        RECT  1.410 -0.165 1.520 0.445 ;
        RECT  0.195 -0.165 1.410 0.165 ;
        RECT  0.085 -0.165 0.195 0.455 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 1.635 1.600 1.965 ;
        RECT  0.575 1.390 0.745 1.965 ;
        RECT  0.195 1.635 0.575 1.965 ;
        RECT  0.085 1.335 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.075 0.255 1.320 0.440 ;
        RECT  0.305 1.210 1.295 1.300 ;
        RECT  0.315 0.275 0.485 0.580 ;
    END
END GAOI22D1

MACRO GBUFFD1
    CLASS CORE ;
    FOREIGN GBUFFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.305 0.750 1.525 ;
        RECT  0.575 0.305 0.650 0.415 ;
        RECT  0.605 1.200 0.650 1.525 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.165 0.800 0.165 ;
        RECT  0.315 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 1.635 0.800 1.965 ;
        RECT  0.315 1.200 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.450 0.510 0.560 0.940 ;
        RECT  0.195 0.510 0.450 0.610 ;
        RECT  0.150 0.265 0.195 0.610 ;
        RECT  0.150 1.200 0.195 1.525 ;
        RECT  0.085 0.265 0.150 1.525 ;
        RECT  0.050 0.510 0.085 1.310 ;
    END
END GBUFFD1

MACRO GBUFFD2
    CLASS CORE ;
    FOREIGN GBUFFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.305 ;
        RECT  1.255 0.510 1.450 0.610 ;
        RECT  1.115 1.205 1.450 1.305 ;
        RECT  1.145 0.275 1.255 0.610 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.095 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  0.995 -0.165 1.375 0.165 ;
        RECT  0.885 -0.165 0.995 0.465 ;
        RECT  0.455 -0.165 0.885 0.165 ;
        RECT  0.345 -0.165 0.455 0.455 ;
        RECT  0.195 -0.165 0.345 0.165 ;
        RECT  0.085 -0.165 0.195 0.455 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.635 1.600 1.965 ;
        RECT  1.375 1.395 1.545 1.965 ;
        RECT  0.995 1.635 1.375 1.965 ;
        RECT  0.885 1.335 0.995 1.965 ;
        RECT  0.195 1.635 0.885 1.965 ;
        RECT  0.195 1.205 0.495 1.315 ;
        RECT  0.085 1.205 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.730 1.360 1.110 ;
        RECT  1.140 1.000 1.250 1.110 ;
        RECT  1.030 0.730 1.140 1.110 ;
        RECT  0.760 1.000 1.030 1.110 ;
        RECT  0.715 0.470 0.760 1.320 ;
        RECT  0.660 0.275 0.715 1.525 ;
        RECT  0.605 0.275 0.660 0.580 ;
        RECT  0.605 1.210 0.660 1.525 ;
        RECT  0.240 0.690 0.350 1.095 ;
    END
END GBUFFD2

MACRO GBUFFD3
    CLASS CORE ;
    FOREIGN GBUFFD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.305 ;
        RECT  1.255 0.510 1.450 0.610 ;
        RECT  0.715 1.205 1.450 1.305 ;
        RECT  1.145 0.275 1.255 0.610 ;
        RECT  0.715 0.510 1.145 0.610 ;
        RECT  0.605 0.275 0.715 0.610 ;
        RECT  0.605 1.205 0.715 1.525 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.510 0.360 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.410 ;
        RECT  0.485 -0.165 0.855 0.165 ;
        RECT  0.315 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.635 1.600 1.965 ;
        RECT  1.375 1.395 1.545 1.965 ;
        RECT  1.025 1.635 1.375 1.965 ;
        RECT  0.855 1.395 1.025 1.965 ;
        RECT  0.485 1.635 0.855 1.965 ;
        RECT  0.315 1.205 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.730 1.360 1.110 ;
        RECT  1.140 1.000 1.250 1.110 ;
        RECT  1.030 0.730 1.140 1.110 ;
        RECT  0.570 1.000 1.030 1.110 ;
        RECT  0.460 0.730 0.570 1.110 ;
        RECT  0.150 1.000 0.460 1.110 ;
        RECT  0.150 0.305 0.225 0.415 ;
        RECT  0.150 1.385 0.225 1.495 ;
        RECT  0.055 0.305 0.150 1.495 ;
    END
END GBUFFD3

MACRO GBUFFD4
    CLASS CORE ;
    FOREIGN GBUFFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 2.350 1.305 ;
        RECT  2.055 0.510 2.250 0.610 ;
        RECT  1.300 1.205 2.250 1.305 ;
        RECT  1.945 0.275 2.055 0.610 ;
        RECT  1.255 0.510 1.945 0.610 ;
        RECT  1.050 1.195 1.300 1.305 ;
        RECT  1.145 0.275 1.255 0.610 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.090 ;
        RECT  0.350 0.980 0.450 1.090 ;
        RECT  0.240 0.690 0.350 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 -0.165 2.400 0.165 ;
        RECT  2.175 -0.165 2.345 0.410 ;
        RECT  1.825 -0.165 2.175 0.165 ;
        RECT  1.655 -0.165 1.825 0.410 ;
        RECT  1.545 -0.165 1.655 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.410 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.635 2.400 1.965 ;
        RECT  2.175 1.395 2.345 1.965 ;
        RECT  1.825 1.635 2.175 1.965 ;
        RECT  1.655 1.395 1.825 1.965 ;
        RECT  1.545 1.635 1.655 1.965 ;
        RECT  1.375 1.395 1.545 1.965 ;
        RECT  1.025 1.635 1.375 1.965 ;
        RECT  0.855 1.395 1.025 1.965 ;
        RECT  0.745 1.635 0.855 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.395 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.050 0.730 2.160 1.110 ;
        RECT  0.955 0.770 2.050 0.880 ;
        RECT  0.845 0.500 0.955 1.305 ;
        RECT  0.455 0.500 0.845 0.600 ;
        RECT  0.315 1.195 0.845 1.305 ;
        RECT  0.345 0.275 0.455 0.600 ;
    END
END GBUFFD4

MACRO GBUFFD8
    CLASS CORE ;
    FOREIGN GBUFFD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.510 4.750 1.305 ;
        RECT  4.455 0.510 4.650 0.610 ;
        RECT  2.100 1.200 4.650 1.305 ;
        RECT  4.345 0.275 4.455 0.610 ;
        RECT  3.655 0.510 4.345 0.610 ;
        RECT  3.545 0.275 3.655 0.610 ;
        RECT  2.855 0.510 3.545 0.610 ;
        RECT  2.745 0.275 2.855 0.610 ;
        RECT  2.055 0.510 2.745 0.610 ;
        RECT  1.850 1.190 2.100 1.305 ;
        RECT  1.945 0.275 2.055 0.610 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.160 1.090 ;
        RECT  0.350 0.770 1.040 0.880 ;
        RECT  0.240 0.690 0.350 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.745 -0.165 4.800 0.165 ;
        RECT  4.575 -0.165 4.745 0.410 ;
        RECT  4.225 -0.165 4.575 0.165 ;
        RECT  4.055 -0.165 4.225 0.410 ;
        RECT  3.945 -0.165 4.055 0.165 ;
        RECT  3.775 -0.165 3.945 0.410 ;
        RECT  3.425 -0.165 3.775 0.165 ;
        RECT  3.255 -0.165 3.425 0.410 ;
        RECT  3.145 -0.165 3.255 0.165 ;
        RECT  2.975 -0.165 3.145 0.410 ;
        RECT  2.625 -0.165 2.975 0.165 ;
        RECT  2.455 -0.165 2.625 0.410 ;
        RECT  2.345 -0.165 2.455 0.165 ;
        RECT  2.175 -0.165 2.345 0.410 ;
        RECT  1.825 -0.165 2.175 0.165 ;
        RECT  1.655 -0.165 1.825 0.410 ;
        RECT  1.545 -0.165 1.655 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.410 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.745 1.635 4.800 1.965 ;
        RECT  4.575 1.395 4.745 1.965 ;
        RECT  4.225 1.635 4.575 1.965 ;
        RECT  4.055 1.395 4.225 1.965 ;
        RECT  3.945 1.635 4.055 1.965 ;
        RECT  3.775 1.395 3.945 1.965 ;
        RECT  3.425 1.635 3.775 1.965 ;
        RECT  3.255 1.395 3.425 1.965 ;
        RECT  3.145 1.635 3.255 1.965 ;
        RECT  2.975 1.395 3.145 1.965 ;
        RECT  2.625 1.635 2.975 1.965 ;
        RECT  2.455 1.395 2.625 1.965 ;
        RECT  2.345 1.635 2.455 1.965 ;
        RECT  2.175 1.395 2.345 1.965 ;
        RECT  1.825 1.635 2.175 1.965 ;
        RECT  1.655 1.395 1.825 1.965 ;
        RECT  1.545 1.635 1.655 1.965 ;
        RECT  1.375 1.395 1.545 1.965 ;
        RECT  1.025 1.635 1.375 1.965 ;
        RECT  0.855 1.395 1.025 1.965 ;
        RECT  0.745 1.635 0.855 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.395 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.450 0.730 4.560 1.110 ;
        RECT  1.755 0.770 4.450 0.880 ;
        RECT  1.645 0.500 1.755 1.305 ;
        RECT  1.255 0.500 1.645 0.600 ;
        RECT  0.315 1.195 1.645 1.305 ;
        RECT  1.250 0.740 1.400 1.090 ;
        RECT  1.145 0.275 1.255 0.600 ;
        RECT  0.455 0.500 1.145 0.600 ;
        RECT  0.345 0.275 0.455 0.600 ;
    END
END GBUFFD8

MACRO GDCAP
    CLASS CORE ;
    FOREIGN GDCAP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 -0.165 0.800 0.165 ;
        RECT  0.345 -0.165 0.455 0.465 ;
        RECT  0.195 -0.165 0.345 0.165 ;
        RECT  0.085 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GDCAP

MACRO GDCAP10
    CLASS CORE ;
    FOREIGN GDCAP10 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.655 -0.165 8.000 0.165 ;
        RECT  7.545 -0.165 7.655 0.465 ;
        RECT  7.395 -0.165 7.545 0.165 ;
        RECT  7.285 -0.165 7.395 0.465 ;
        RECT  6.855 -0.165 7.285 0.165 ;
        RECT  6.745 -0.165 6.855 0.465 ;
        RECT  6.595 -0.165 6.745 0.165 ;
        RECT  6.485 -0.165 6.595 0.465 ;
        RECT  6.055 -0.165 6.485 0.165 ;
        RECT  5.945 -0.165 6.055 0.465 ;
        RECT  5.795 -0.165 5.945 0.165 ;
        RECT  5.685 -0.165 5.795 0.465 ;
        RECT  5.255 -0.165 5.685 0.165 ;
        RECT  5.145 -0.165 5.255 0.465 ;
        RECT  4.995 -0.165 5.145 0.165 ;
        RECT  4.885 -0.165 4.995 0.465 ;
        RECT  4.455 -0.165 4.885 0.165 ;
        RECT  4.345 -0.165 4.455 0.465 ;
        RECT  4.195 -0.165 4.345 0.165 ;
        RECT  4.085 -0.165 4.195 0.465 ;
        RECT  3.655 -0.165 4.085 0.165 ;
        RECT  3.545 -0.165 3.655 0.465 ;
        RECT  3.395 -0.165 3.545 0.165 ;
        RECT  3.285 -0.165 3.395 0.465 ;
        RECT  2.855 -0.165 3.285 0.165 ;
        RECT  2.745 -0.165 2.855 0.465 ;
        RECT  2.595 -0.165 2.745 0.165 ;
        RECT  2.485 -0.165 2.595 0.465 ;
        RECT  2.055 -0.165 2.485 0.165 ;
        RECT  1.945 -0.165 2.055 0.465 ;
        RECT  1.795 -0.165 1.945 0.165 ;
        RECT  1.685 -0.165 1.795 0.465 ;
        RECT  1.255 -0.165 1.685 0.165 ;
        RECT  1.145 -0.165 1.255 0.465 ;
        RECT  0.995 -0.165 1.145 0.165 ;
        RECT  0.885 -0.165 0.995 0.465 ;
        RECT  0.455 -0.165 0.885 0.165 ;
        RECT  0.345 -0.165 0.455 0.465 ;
        RECT  0.195 -0.165 0.345 0.165 ;
        RECT  0.085 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.915 1.635 8.000 1.965 ;
        RECT  7.805 1.200 7.915 1.965 ;
        RECT  7.505 1.200 7.805 1.310 ;
        RECT  7.115 1.635 7.805 1.965 ;
        RECT  7.005 1.200 7.115 1.965 ;
        RECT  6.705 1.200 7.005 1.310 ;
        RECT  6.315 1.635 7.005 1.965 ;
        RECT  6.205 1.200 6.315 1.965 ;
        RECT  5.905 1.200 6.205 1.310 ;
        RECT  5.515 1.635 6.205 1.965 ;
        RECT  5.405 1.200 5.515 1.965 ;
        RECT  5.105 1.200 5.405 1.310 ;
        RECT  4.715 1.635 5.405 1.965 ;
        RECT  4.605 1.200 4.715 1.965 ;
        RECT  4.305 1.200 4.605 1.310 ;
        RECT  3.915 1.635 4.605 1.965 ;
        RECT  3.805 1.200 3.915 1.965 ;
        RECT  3.505 1.200 3.805 1.310 ;
        RECT  3.115 1.635 3.805 1.965 ;
        RECT  3.005 1.200 3.115 1.965 ;
        RECT  2.705 1.200 3.005 1.310 ;
        RECT  2.315 1.635 3.005 1.965 ;
        RECT  2.205 1.200 2.315 1.965 ;
        RECT  1.905 1.200 2.205 1.310 ;
        RECT  1.515 1.635 2.205 1.965 ;
        RECT  1.405 1.200 1.515 1.965 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  0.715 1.635 1.405 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.805 0.275 7.915 0.650 ;
        RECT  7.540 0.560 7.805 0.650 ;
        RECT  7.660 0.740 7.770 1.110 ;
        RECT  7.395 1.020 7.660 1.110 ;
        RECT  7.430 0.560 7.540 0.910 ;
        RECT  7.115 0.560 7.430 0.650 ;
        RECT  7.285 1.020 7.395 1.525 ;
        RECT  6.970 1.020 7.285 1.110 ;
        RECT  7.005 0.275 7.115 0.650 ;
        RECT  6.740 0.560 7.005 0.650 ;
        RECT  6.860 0.740 6.970 1.110 ;
        RECT  6.595 1.020 6.860 1.110 ;
        RECT  6.630 0.560 6.740 0.910 ;
        RECT  6.315 0.560 6.630 0.650 ;
        RECT  6.485 1.020 6.595 1.525 ;
        RECT  6.170 1.020 6.485 1.110 ;
        RECT  6.205 0.275 6.315 0.650 ;
        RECT  5.940 0.560 6.205 0.650 ;
        RECT  6.060 0.740 6.170 1.110 ;
        RECT  5.795 1.020 6.060 1.110 ;
        RECT  5.830 0.560 5.940 0.910 ;
        RECT  5.515 0.560 5.830 0.650 ;
        RECT  5.685 1.020 5.795 1.525 ;
        RECT  5.370 1.020 5.685 1.110 ;
        RECT  5.405 0.275 5.515 0.650 ;
        RECT  5.140 0.560 5.405 0.650 ;
        RECT  5.260 0.740 5.370 1.110 ;
        RECT  4.995 1.020 5.260 1.110 ;
        RECT  5.030 0.560 5.140 0.910 ;
        RECT  4.715 0.560 5.030 0.650 ;
        RECT  4.885 1.020 4.995 1.525 ;
        RECT  4.570 1.020 4.885 1.110 ;
        RECT  4.605 0.275 4.715 0.650 ;
        RECT  4.340 0.560 4.605 0.650 ;
        RECT  4.460 0.740 4.570 1.110 ;
        RECT  4.195 1.020 4.460 1.110 ;
        RECT  4.230 0.560 4.340 0.910 ;
        RECT  3.915 0.560 4.230 0.650 ;
        RECT  4.085 1.020 4.195 1.525 ;
        RECT  3.770 1.020 4.085 1.110 ;
        RECT  3.805 0.275 3.915 0.650 ;
        RECT  3.540 0.560 3.805 0.650 ;
        RECT  3.660 0.740 3.770 1.110 ;
        RECT  3.395 1.020 3.660 1.110 ;
        RECT  3.430 0.560 3.540 0.910 ;
        RECT  3.115 0.560 3.430 0.650 ;
        RECT  3.285 1.020 3.395 1.525 ;
        RECT  2.970 1.020 3.285 1.110 ;
        RECT  3.005 0.275 3.115 0.650 ;
        RECT  2.740 0.560 3.005 0.650 ;
        RECT  2.860 0.740 2.970 1.110 ;
        RECT  2.595 1.020 2.860 1.110 ;
        RECT  2.630 0.560 2.740 0.910 ;
        RECT  2.315 0.560 2.630 0.650 ;
        RECT  2.485 1.020 2.595 1.525 ;
        RECT  2.170 1.020 2.485 1.110 ;
        RECT  2.205 0.275 2.315 0.650 ;
        RECT  1.940 0.560 2.205 0.650 ;
        RECT  2.060 0.740 2.170 1.110 ;
        RECT  1.795 1.020 2.060 1.110 ;
        RECT  1.830 0.560 1.940 0.910 ;
        RECT  1.515 0.560 1.830 0.650 ;
        RECT  1.685 1.020 1.795 1.525 ;
        RECT  1.370 1.020 1.685 1.110 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GDCAP10

MACRO GDCAP2
    CLASS CORE ;
    FOREIGN GDCAP2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.255 -0.165 1.600 0.165 ;
        RECT  1.145 -0.165 1.255 0.465 ;
        RECT  0.995 -0.165 1.145 0.165 ;
        RECT  0.885 -0.165 0.995 0.465 ;
        RECT  0.455 -0.165 0.885 0.165 ;
        RECT  0.345 -0.165 0.455 0.465 ;
        RECT  0.195 -0.165 0.345 0.165 ;
        RECT  0.085 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.200 1.515 1.965 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  0.715 1.635 1.405 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GDCAP2

MACRO GDCAP3
    CLASS CORE ;
    FOREIGN GDCAP3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 -0.165 2.400 0.165 ;
        RECT  1.945 -0.165 2.055 0.465 ;
        RECT  1.795 -0.165 1.945 0.165 ;
        RECT  1.685 -0.165 1.795 0.465 ;
        RECT  1.255 -0.165 1.685 0.165 ;
        RECT  1.145 -0.165 1.255 0.465 ;
        RECT  0.995 -0.165 1.145 0.165 ;
        RECT  0.885 -0.165 0.995 0.465 ;
        RECT  0.455 -0.165 0.885 0.165 ;
        RECT  0.345 -0.165 0.455 0.465 ;
        RECT  0.195 -0.165 0.345 0.165 ;
        RECT  0.085 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 1.635 2.400 1.965 ;
        RECT  2.205 1.200 2.315 1.965 ;
        RECT  1.905 1.200 2.205 1.310 ;
        RECT  1.515 1.635 2.205 1.965 ;
        RECT  1.405 1.200 1.515 1.965 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  0.715 1.635 1.405 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.275 2.315 0.650 ;
        RECT  1.940 0.560 2.205 0.650 ;
        RECT  2.060 0.740 2.170 1.110 ;
        RECT  1.795 1.020 2.060 1.110 ;
        RECT  1.830 0.560 1.940 0.910 ;
        RECT  1.515 0.560 1.830 0.650 ;
        RECT  1.685 1.020 1.795 1.525 ;
        RECT  1.370 1.020 1.685 1.110 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GDCAP3

MACRO GDCAP4
    CLASS CORE ;
    FOREIGN GDCAP4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.855 -0.165 3.200 0.165 ;
        RECT  2.745 -0.165 2.855 0.465 ;
        RECT  2.595 -0.165 2.745 0.165 ;
        RECT  2.485 -0.165 2.595 0.465 ;
        RECT  2.055 -0.165 2.485 0.165 ;
        RECT  1.945 -0.165 2.055 0.465 ;
        RECT  1.795 -0.165 1.945 0.165 ;
        RECT  1.685 -0.165 1.795 0.465 ;
        RECT  1.255 -0.165 1.685 0.165 ;
        RECT  1.145 -0.165 1.255 0.465 ;
        RECT  0.995 -0.165 1.145 0.165 ;
        RECT  0.885 -0.165 0.995 0.465 ;
        RECT  0.455 -0.165 0.885 0.165 ;
        RECT  0.345 -0.165 0.455 0.465 ;
        RECT  0.195 -0.165 0.345 0.165 ;
        RECT  0.085 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.115 1.635 3.200 1.965 ;
        RECT  3.005 1.200 3.115 1.965 ;
        RECT  2.705 1.200 3.005 1.310 ;
        RECT  2.315 1.635 3.005 1.965 ;
        RECT  2.205 1.200 2.315 1.965 ;
        RECT  1.905 1.200 2.205 1.310 ;
        RECT  1.515 1.635 2.205 1.965 ;
        RECT  1.405 1.200 1.515 1.965 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  0.715 1.635 1.405 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.005 0.275 3.115 0.650 ;
        RECT  2.740 0.560 3.005 0.650 ;
        RECT  2.860 0.740 2.970 1.110 ;
        RECT  2.595 1.020 2.860 1.110 ;
        RECT  2.630 0.560 2.740 0.910 ;
        RECT  2.315 0.560 2.630 0.650 ;
        RECT  2.485 1.020 2.595 1.525 ;
        RECT  2.170 1.020 2.485 1.110 ;
        RECT  2.205 0.275 2.315 0.650 ;
        RECT  1.940 0.560 2.205 0.650 ;
        RECT  2.060 0.740 2.170 1.110 ;
        RECT  1.795 1.020 2.060 1.110 ;
        RECT  1.830 0.560 1.940 0.910 ;
        RECT  1.515 0.560 1.830 0.650 ;
        RECT  1.685 1.020 1.795 1.525 ;
        RECT  1.370 1.020 1.685 1.110 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GDCAP4

MACRO GDFCNQD1
    CLASS CORE ;
    FOREIGN GDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.305 5.550 1.495 ;
        RECT  5.375 0.305 5.450 0.415 ;
        RECT  5.375 1.385 5.450 1.495 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.755 0.910 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.540 2.960 0.910 ;
        RECT  1.500 0.540 2.850 0.630 ;
        RECT  1.410 0.540 1.500 0.680 ;
        RECT  1.370 0.590 1.410 0.680 ;
        RECT  1.260 0.590 1.370 0.920 ;
        RECT  0.955 0.590 1.260 0.680 ;
        RECT  0.865 0.510 0.955 0.680 ;
        RECT  0.355 0.510 0.865 0.600 ;
        RECT  0.240 0.510 0.355 0.910 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.420 0.600 4.580 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.265 -0.165 5.600 0.165 ;
        RECT  5.135 -0.165 5.265 0.495 ;
        RECT  4.190 -0.165 5.135 0.165 ;
        RECT  4.080 -0.165 4.190 0.445 ;
        RECT  2.865 -0.165 4.080 0.165 ;
        RECT  2.735 -0.165 2.865 0.445 ;
        RECT  2.330 -0.165 2.735 0.165 ;
        RECT  2.215 -0.165 2.330 0.450 ;
        RECT  0.485 -0.165 2.215 0.165 ;
        RECT  0.315 -0.165 0.485 0.415 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.635 5.600 1.965 ;
        RECT  5.135 1.150 5.270 1.965 ;
        RECT  4.485 1.635 5.135 1.965 ;
        RECT  4.315 1.210 4.485 1.965 ;
        RECT  2.885 1.635 4.315 1.965 ;
        RECT  2.715 1.210 2.885 1.965 ;
        RECT  2.085 1.635 2.715 1.965 ;
        RECT  1.915 1.210 2.085 1.965 ;
        RECT  0.485 1.635 1.915 1.965 ;
        RECT  0.315 1.210 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.760 0.740 5.360 0.910 ;
        RECT  4.850 1.210 5.030 1.525 ;
        RECT  4.850 0.255 5.015 0.630 ;
        RECT  4.670 0.295 4.760 1.525 ;
        RECT  4.575 0.295 4.670 0.420 ;
        RECT  4.580 1.210 4.670 1.525 ;
        RECT  4.305 0.255 4.485 0.490 ;
        RECT  4.035 0.740 4.330 0.910 ;
        RECT  4.035 1.215 4.215 1.525 ;
        RECT  3.945 0.540 4.035 1.110 ;
        RECT  3.745 0.255 3.990 0.450 ;
        RECT  3.655 0.540 3.945 0.630 ;
        RECT  3.655 1.010 3.945 1.110 ;
        RECT  3.780 1.210 3.925 1.525 ;
        RECT  3.620 0.720 3.840 0.920 ;
        RECT  3.545 0.275 3.655 0.630 ;
        RECT  3.545 1.010 3.655 1.360 ;
        RECT  3.150 0.740 3.530 0.910 ;
        RECT  3.250 0.255 3.435 0.650 ;
        RECT  3.250 1.210 3.420 1.510 ;
        RECT  3.050 0.300 3.150 1.505 ;
        RECT  2.975 0.300 3.050 0.425 ;
        RECT  2.975 1.380 3.050 1.505 ;
        RECT  2.630 0.730 2.740 1.110 ;
        RECT  2.420 0.255 2.645 0.450 ;
        RECT  1.255 1.010 2.630 1.110 ;
        RECT  2.450 1.210 2.620 1.510 ;
        RECT  2.175 1.210 2.355 1.510 ;
        RECT  2.050 0.730 2.350 0.910 ;
        RECT  1.905 0.255 2.125 0.450 ;
        RECT  1.715 0.740 1.950 0.920 ;
        RECT  1.645 1.210 1.825 1.510 ;
        RECT  1.410 0.275 1.815 0.445 ;
        RECT  1.365 1.210 1.545 1.510 ;
        RECT  1.115 0.255 1.320 0.500 ;
        RECT  1.145 1.010 1.255 1.350 ;
        RECT  0.955 0.770 1.170 0.880 ;
        RECT  0.850 1.210 1.030 1.510 ;
        RECT  0.575 0.305 1.025 0.415 ;
        RECT  0.865 0.770 0.955 1.110 ;
        RECT  0.145 1.020 0.865 1.110 ;
        RECT  0.575 1.210 0.755 1.510 ;
        RECT  0.145 0.305 0.225 0.415 ;
        RECT  0.145 1.385 0.225 1.495 ;
        RECT  0.050 0.305 0.145 1.495 ;
        LAYER VIA1 ;
        RECT  4.890 1.210 4.990 1.310 ;
        RECT  4.850 0.390 4.950 0.490 ;
        RECT  4.620 1.410 4.720 1.510 ;
        RECT  4.450 0.950 4.550 1.050 ;
        RECT  4.075 1.410 4.175 1.510 ;
        RECT  3.820 0.340 3.920 0.440 ;
        RECT  3.815 1.250 3.915 1.350 ;
        RECT  3.695 0.750 3.795 0.850 ;
        RECT  3.290 0.550 3.390 0.650 ;
        RECT  3.250 1.250 3.350 1.350 ;
        RECT  2.850 0.710 2.950 0.810 ;
        RECT  2.480 1.250 2.580 1.350 ;
        RECT  2.470 0.340 2.570 0.440 ;
        RECT  2.250 0.770 2.350 0.870 ;
        RECT  2.215 1.410 2.315 1.510 ;
        RECT  1.850 0.780 1.950 0.880 ;
        RECT  1.685 1.410 1.785 1.510 ;
        RECT  1.405 1.210 1.505 1.310 ;
        RECT  1.290 1.010 1.390 1.110 ;
        RECT  1.175 0.310 1.275 0.410 ;
        RECT  0.890 1.410 0.990 1.510 ;
        RECT  0.650 1.250 0.750 1.350 ;
        LAYER M2 ;
        RECT  4.950 1.210 5.030 1.310 ;
        RECT  4.850 0.350 4.950 1.310 ;
        RECT  4.250 0.350 4.850 0.450 ;
        RECT  3.915 1.210 4.850 1.310 ;
        RECT  4.035 1.410 4.760 1.510 ;
        RECT  4.450 0.910 4.550 1.110 ;
        RECT  2.350 1.010 4.450 1.110 ;
        RECT  4.150 0.350 4.250 0.650 ;
        RECT  3.250 0.550 4.150 0.650 ;
        RECT  1.950 0.340 3.960 0.440 ;
        RECT  3.815 1.210 3.915 1.390 ;
        RECT  2.950 0.750 3.835 0.850 ;
        RECT  3.250 1.210 3.350 1.390 ;
        RECT  2.580 1.210 3.250 1.310 ;
        RECT  2.850 0.670 2.950 0.850 ;
        RECT  2.480 1.210 2.580 1.390 ;
        RECT  1.950 1.210 2.480 1.310 ;
        RECT  0.850 1.410 2.355 1.510 ;
        RECT  2.250 0.730 2.350 1.110 ;
        RECT  1.850 0.340 1.950 1.310 ;
        RECT  1.135 1.210 1.545 1.310 ;
        RECT  1.350 1.010 1.430 1.110 ;
        RECT  1.250 0.310 1.350 1.110 ;
        RECT  1.135 0.310 1.250 0.410 ;
        RECT  1.035 1.110 1.135 1.310 ;
        RECT  0.750 1.110 1.035 1.210 ;
        RECT  0.650 1.110 0.750 1.390 ;
    END
END GDFCNQD1

MACRO GDFQD1
    CLASS CORE ;
    FOREIGN GDFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.305 4.750 1.495 ;
        RECT  4.575 0.305 4.650 0.415 ;
        RECT  4.575 1.385 4.650 1.495 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.755 0.910 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.740 3.550 1.090 ;
        RECT  2.770 1.000 3.440 1.090 ;
        RECT  2.680 0.770 2.770 1.090 ;
        RECT  2.545 0.770 2.680 0.880 ;
        RECT  2.455 0.540 2.545 0.880 ;
        RECT  1.705 0.540 2.455 0.630 ;
        RECT  1.615 0.540 1.705 0.680 ;
        RECT  1.370 0.590 1.615 0.680 ;
        RECT  1.260 0.590 1.370 0.920 ;
        RECT  0.955 0.590 1.260 0.680 ;
        RECT  0.865 0.510 0.955 0.680 ;
        RECT  0.355 0.510 0.865 0.600 ;
        RECT  0.240 0.510 0.355 0.910 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.455 -0.165 4.800 0.165 ;
        RECT  4.345 -0.165 4.455 0.445 ;
        RECT  3.655 -0.165 4.345 0.165 ;
        RECT  3.545 -0.165 3.655 0.445 ;
        RECT  2.055 -0.165 3.545 0.165 ;
        RECT  1.945 -0.165 2.055 0.445 ;
        RECT  0.485 -0.165 1.945 0.165 ;
        RECT  0.315 -0.165 0.485 0.415 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.485 1.635 4.800 1.965 ;
        RECT  4.315 1.210 4.485 1.965 ;
        RECT  3.685 1.635 4.315 1.965 ;
        RECT  3.515 1.210 3.685 1.965 ;
        RECT  2.055 1.635 3.515 1.965 ;
        RECT  2.055 1.210 2.085 1.320 ;
        RECT  1.945 1.210 2.055 1.965 ;
        RECT  1.915 1.210 1.945 1.320 ;
        RECT  0.485 1.635 1.945 1.965 ;
        RECT  0.315 1.210 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.470 0.560 4.560 1.090 ;
        RECT  4.195 0.560 4.470 0.650 ;
        RECT  4.195 1.000 4.470 1.090 ;
        RECT  3.980 0.770 4.380 0.880 ;
        RECT  4.085 0.275 4.195 0.650 ;
        RECT  4.085 1.000 4.195 1.525 ;
        RECT  3.770 1.000 4.085 1.090 ;
        RECT  3.745 0.265 3.995 0.445 ;
        RECT  3.890 0.535 3.980 0.880 ;
        RECT  3.805 1.210 3.950 1.525 ;
        RECT  3.475 0.535 3.890 0.645 ;
        RECT  3.660 0.740 3.770 1.090 ;
        RECT  3.250 1.210 3.405 1.525 ;
        RECT  3.350 0.275 3.395 0.445 ;
        RECT  3.260 0.275 3.350 0.910 ;
        RECT  2.860 0.740 3.260 0.910 ;
        RECT  2.975 0.255 3.155 0.500 ;
        RECT  3.010 1.180 3.150 1.525 ;
        RECT  2.710 1.180 2.890 1.525 ;
        RECT  2.715 0.275 2.885 0.640 ;
        RECT  2.705 0.540 2.715 0.640 ;
        RECT  2.350 0.305 2.625 0.415 ;
        RECT  2.450 1.100 2.590 1.525 ;
        RECT  2.175 0.265 2.350 0.445 ;
        RECT  2.195 1.220 2.350 1.525 ;
        RECT  2.060 0.730 2.170 1.110 ;
        RECT  1.255 1.010 2.060 1.110 ;
        RECT  1.830 0.730 1.950 0.920 ;
        RECT  1.640 0.800 1.830 0.920 ;
        RECT  1.515 0.305 1.825 0.415 ;
        RECT  1.645 1.210 1.825 1.510 ;
        RECT  1.365 1.210 1.545 1.510 ;
        RECT  1.405 0.275 1.515 0.445 ;
        RECT  1.135 0.255 1.315 0.500 ;
        RECT  1.145 1.010 1.255 1.350 ;
        RECT  0.955 0.770 1.170 0.880 ;
        RECT  1.110 1.010 1.145 1.110 ;
        RECT  0.850 1.210 1.030 1.510 ;
        RECT  0.575 0.305 1.025 0.415 ;
        RECT  0.865 0.770 0.955 1.110 ;
        RECT  0.145 1.020 0.865 1.110 ;
        RECT  0.575 1.210 0.755 1.490 ;
        RECT  0.145 0.305 0.225 0.415 ;
        RECT  0.145 1.385 0.225 1.495 ;
        RECT  0.055 0.305 0.145 1.495 ;
        LAYER VIA1 ;
        RECT  3.850 1.350 3.950 1.450 ;
        RECT  3.810 0.300 3.910 0.400 ;
        RECT  3.515 0.540 3.615 0.640 ;
        RECT  3.250 1.370 3.350 1.470 ;
        RECT  3.210 0.775 3.310 0.875 ;
        RECT  3.050 1.220 3.150 1.320 ;
        RECT  3.015 0.300 3.115 0.400 ;
        RECT  2.750 1.205 2.850 1.305 ;
        RECT  2.745 0.540 2.845 0.640 ;
        RECT  2.450 1.140 2.550 1.240 ;
        RECT  2.250 0.305 2.350 0.405 ;
        RECT  2.250 1.350 2.350 1.450 ;
        RECT  1.810 0.820 1.910 0.920 ;
        RECT  1.685 1.410 1.785 1.510 ;
        RECT  1.405 1.210 1.505 1.310 ;
        RECT  1.175 0.310 1.275 0.410 ;
        RECT  1.150 1.010 1.250 1.110 ;
        RECT  0.890 1.410 0.990 1.510 ;
        RECT  0.615 1.210 0.715 1.310 ;
        LAYER M2 ;
        RECT  3.850 0.300 3.950 1.490 ;
        RECT  2.550 0.300 3.850 0.400 ;
        RECT  2.860 0.540 3.655 0.640 ;
        RECT  3.250 0.775 3.350 1.510 ;
        RECT  3.170 0.775 3.250 0.875 ;
        RECT  3.050 1.180 3.150 1.510 ;
        RECT  2.350 1.410 3.050 1.510 ;
        RECT  2.860 1.205 2.890 1.305 ;
        RECT  2.760 0.540 2.860 1.305 ;
        RECT  2.705 0.540 2.760 0.640 ;
        RECT  2.710 1.205 2.760 1.305 ;
        RECT  2.450 0.300 2.550 1.280 ;
        RECT  2.250 0.265 2.350 1.510 ;
        RECT  1.770 0.820 2.250 0.920 ;
        RECT  0.850 1.410 1.825 1.510 ;
        RECT  0.575 1.210 1.545 1.310 ;
        RECT  1.250 0.310 1.350 1.110 ;
        RECT  1.135 0.310 1.250 0.410 ;
        RECT  1.110 1.010 1.250 1.110 ;
    END
END GDFQD1

MACRO GFILL
    CLASS CORE ;
    FOREIGN GFILL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 0.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 0.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.605 1.200 0.715 1.525 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.085 0.275 0.485 0.465 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GFILL

MACRO GFILL10
    CLASS CORE ;
    FOREIGN GFILL10 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 8.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 8.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.805 0.275 7.915 0.650 ;
        RECT  7.805 1.200 7.915 1.525 ;
        RECT  7.540 0.560 7.805 0.650 ;
        RECT  7.505 1.200 7.805 1.310 ;
        RECT  7.660 0.740 7.770 1.110 ;
        RECT  7.285 0.275 7.685 0.465 ;
        RECT  7.395 1.020 7.660 1.110 ;
        RECT  7.430 0.560 7.540 0.910 ;
        RECT  7.115 0.560 7.430 0.650 ;
        RECT  7.285 1.020 7.395 1.525 ;
        RECT  6.970 1.020 7.285 1.110 ;
        RECT  7.005 0.275 7.115 0.650 ;
        RECT  7.005 1.200 7.115 1.525 ;
        RECT  6.740 0.560 7.005 0.650 ;
        RECT  6.705 1.200 7.005 1.310 ;
        RECT  6.860 0.740 6.970 1.110 ;
        RECT  6.485 0.275 6.885 0.465 ;
        RECT  6.595 1.020 6.860 1.110 ;
        RECT  6.630 0.560 6.740 0.910 ;
        RECT  6.315 0.560 6.630 0.650 ;
        RECT  6.485 1.020 6.595 1.525 ;
        RECT  6.170 1.020 6.485 1.110 ;
        RECT  6.205 0.275 6.315 0.650 ;
        RECT  6.205 1.200 6.315 1.525 ;
        RECT  5.940 0.560 6.205 0.650 ;
        RECT  5.905 1.200 6.205 1.310 ;
        RECT  6.060 0.740 6.170 1.110 ;
        RECT  5.685 0.275 6.085 0.465 ;
        RECT  5.795 1.020 6.060 1.110 ;
        RECT  5.830 0.560 5.940 0.910 ;
        RECT  5.515 0.560 5.830 0.650 ;
        RECT  5.685 1.020 5.795 1.525 ;
        RECT  5.370 1.020 5.685 1.110 ;
        RECT  5.405 0.275 5.515 0.650 ;
        RECT  5.405 1.200 5.515 1.525 ;
        RECT  5.140 0.560 5.405 0.650 ;
        RECT  5.105 1.200 5.405 1.310 ;
        RECT  5.260 0.740 5.370 1.110 ;
        RECT  4.885 0.275 5.285 0.465 ;
        RECT  4.995 1.020 5.260 1.110 ;
        RECT  5.030 0.560 5.140 0.910 ;
        RECT  4.715 0.560 5.030 0.650 ;
        RECT  4.885 1.020 4.995 1.525 ;
        RECT  4.570 1.020 4.885 1.110 ;
        RECT  4.605 0.275 4.715 0.650 ;
        RECT  4.605 1.200 4.715 1.525 ;
        RECT  4.340 0.560 4.605 0.650 ;
        RECT  4.305 1.200 4.605 1.310 ;
        RECT  4.460 0.740 4.570 1.110 ;
        RECT  4.085 0.275 4.485 0.465 ;
        RECT  4.195 1.020 4.460 1.110 ;
        RECT  4.230 0.560 4.340 0.910 ;
        RECT  3.915 0.560 4.230 0.650 ;
        RECT  4.085 1.020 4.195 1.525 ;
        RECT  3.770 1.020 4.085 1.110 ;
        RECT  3.805 0.275 3.915 0.650 ;
        RECT  3.805 1.200 3.915 1.525 ;
        RECT  3.540 0.560 3.805 0.650 ;
        RECT  3.505 1.200 3.805 1.310 ;
        RECT  3.660 0.740 3.770 1.110 ;
        RECT  3.285 0.275 3.685 0.465 ;
        RECT  3.395 1.020 3.660 1.110 ;
        RECT  3.430 0.560 3.540 0.910 ;
        RECT  3.115 0.560 3.430 0.650 ;
        RECT  3.285 1.020 3.395 1.525 ;
        RECT  2.970 1.020 3.285 1.110 ;
        RECT  3.005 0.275 3.115 0.650 ;
        RECT  3.005 1.200 3.115 1.525 ;
        RECT  2.740 0.560 3.005 0.650 ;
        RECT  2.705 1.200 3.005 1.310 ;
        RECT  2.860 0.740 2.970 1.110 ;
        RECT  2.485 0.275 2.885 0.465 ;
        RECT  2.595 1.020 2.860 1.110 ;
        RECT  2.630 0.560 2.740 0.910 ;
        RECT  2.315 0.560 2.630 0.650 ;
        RECT  2.485 1.020 2.595 1.525 ;
        RECT  2.170 1.020 2.485 1.110 ;
        RECT  2.205 0.275 2.315 0.650 ;
        RECT  2.205 1.200 2.315 1.525 ;
        RECT  1.940 0.560 2.205 0.650 ;
        RECT  1.905 1.200 2.205 1.310 ;
        RECT  2.060 0.740 2.170 1.110 ;
        RECT  1.685 0.275 2.085 0.465 ;
        RECT  1.795 1.020 2.060 1.110 ;
        RECT  1.830 0.560 1.940 0.910 ;
        RECT  1.515 0.560 1.830 0.650 ;
        RECT  1.685 1.020 1.795 1.525 ;
        RECT  1.370 1.020 1.685 1.110 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.405 1.200 1.515 1.525 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.885 0.275 1.285 0.465 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.605 1.200 0.715 1.525 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.085 0.275 0.485 0.465 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GFILL10

MACRO GFILL2
    CLASS CORE ;
    FOREIGN GFILL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.405 1.200 1.515 1.525 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.885 0.275 1.285 0.465 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.605 1.200 0.715 1.525 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.085 0.275 0.485 0.465 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GFILL2

MACRO GFILL3
    CLASS CORE ;
    FOREIGN GFILL3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.275 2.315 0.650 ;
        RECT  2.205 1.200 2.315 1.525 ;
        RECT  1.940 0.560 2.205 0.650 ;
        RECT  1.905 1.200 2.205 1.310 ;
        RECT  2.060 0.740 2.170 1.110 ;
        RECT  1.685 0.275 2.085 0.465 ;
        RECT  1.795 1.020 2.060 1.110 ;
        RECT  1.830 0.560 1.940 0.910 ;
        RECT  1.515 0.560 1.830 0.650 ;
        RECT  1.685 1.020 1.795 1.525 ;
        RECT  1.370 1.020 1.685 1.110 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.405 1.200 1.515 1.525 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.885 0.275 1.285 0.465 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.605 1.200 0.715 1.525 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.085 0.275 0.485 0.465 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GFILL3

MACRO GFILL4
    CLASS CORE ;
    FOREIGN GFILL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.200 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.005 0.275 3.115 0.650 ;
        RECT  3.005 1.200 3.115 1.525 ;
        RECT  2.740 0.560 3.005 0.650 ;
        RECT  2.705 1.200 3.005 1.310 ;
        RECT  2.860 0.740 2.970 1.110 ;
        RECT  2.485 0.275 2.885 0.465 ;
        RECT  2.595 1.020 2.860 1.110 ;
        RECT  2.630 0.560 2.740 0.910 ;
        RECT  2.315 0.560 2.630 0.650 ;
        RECT  2.485 1.020 2.595 1.525 ;
        RECT  2.170 1.020 2.485 1.110 ;
        RECT  2.205 0.275 2.315 0.650 ;
        RECT  2.205 1.200 2.315 1.525 ;
        RECT  1.940 0.560 2.205 0.650 ;
        RECT  1.905 1.200 2.205 1.310 ;
        RECT  2.060 0.740 2.170 1.110 ;
        RECT  1.685 0.275 2.085 0.465 ;
        RECT  1.795 1.020 2.060 1.110 ;
        RECT  1.830 0.560 1.940 0.910 ;
        RECT  1.515 0.560 1.830 0.650 ;
        RECT  1.685 1.020 1.795 1.525 ;
        RECT  1.370 1.020 1.685 1.110 ;
        RECT  1.405 0.275 1.515 0.650 ;
        RECT  1.405 1.200 1.515 1.525 ;
        RECT  1.140 0.560 1.405 0.650 ;
        RECT  1.105 1.200 1.405 1.310 ;
        RECT  1.260 0.740 1.370 1.110 ;
        RECT  0.885 0.275 1.285 0.465 ;
        RECT  0.995 1.020 1.260 1.110 ;
        RECT  1.030 0.560 1.140 0.910 ;
        RECT  0.715 0.560 1.030 0.650 ;
        RECT  0.885 1.020 0.995 1.525 ;
        RECT  0.570 1.020 0.885 1.110 ;
        RECT  0.605 0.275 0.715 0.650 ;
        RECT  0.605 1.200 0.715 1.525 ;
        RECT  0.340 0.560 0.605 0.650 ;
        RECT  0.305 1.200 0.605 1.310 ;
        RECT  0.460 0.740 0.570 1.110 ;
        RECT  0.085 0.275 0.485 0.465 ;
        RECT  0.195 1.020 0.460 1.110 ;
        RECT  0.230 0.560 0.340 0.910 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GFILL4

MACRO GINVD1
    CLASS CORE ;
    FOREIGN GINVD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.265 0.195 0.610 ;
        RECT  0.150 1.200 0.195 1.525 ;
        RECT  0.085 0.265 0.150 1.525 ;
        RECT  0.050 0.510 0.085 1.525 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 0.800 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.485 -0.165 0.575 0.165 ;
        RECT  0.315 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.315 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.450 0.710 0.570 1.090 ;
    END
END GINVD1

MACRO GINVD2
    CLASS CORE ;
    FOREIGN GINVD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.190 0.550 1.305 ;
        RECT  0.345 0.275 0.455 0.610 ;
        RECT  0.150 0.510 0.345 0.610 ;
        RECT  0.050 0.510 0.150 1.305 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 0.770 0.640 0.880 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 0.800 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 1.635 0.800 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.395 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
END GINVD2

MACRO GINVD3
    CLASS CORE ;
    FOREIGN GINVD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.305 1.025 0.415 ;
        RECT  0.885 1.200 0.995 1.525 ;
        RECT  0.840 0.305 0.950 0.610 ;
        RECT  0.150 1.200 0.885 1.305 ;
        RECT  0.455 0.510 0.840 0.610 ;
        RECT  0.345 0.275 0.455 0.610 ;
        RECT  0.150 0.510 0.345 0.610 ;
        RECT  0.050 0.510 0.150 1.305 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.160 1.090 ;
        RECT  0.360 0.770 1.040 0.880 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.285 -0.165 1.375 0.165 ;
        RECT  1.115 -0.165 1.285 0.410 ;
        RECT  0.745 -0.165 1.115 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.200 1.515 1.965 ;
        RECT  1.115 1.200 1.405 1.310 ;
        RECT  0.745 1.635 1.405 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.395 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.740 1.400 1.090 ;
    END
END GINVD3

MACRO GINVD4
    CLASS CORE ;
    FOREIGN GINVD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.200 1.295 1.305 ;
        RECT  1.145 0.275 1.255 0.610 ;
        RECT  0.455 0.510 1.145 0.610 ;
        RECT  0.345 0.275 0.455 0.610 ;
        RECT  0.150 0.510 0.345 0.610 ;
        RECT  0.050 0.510 0.150 1.305 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 0.770 1.440 0.880 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.410 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.355 1.515 1.965 ;
        RECT  1.025 1.635 1.405 1.965 ;
        RECT  0.855 1.395 1.025 1.965 ;
        RECT  0.745 1.635 0.855 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.395 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
END GINVD4

MACRO GINVD8
    CLASS CORE ;
    FOREIGN GINVD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.200 2.895 1.305 ;
        RECT  2.745 0.275 2.855 0.610 ;
        RECT  2.055 0.510 2.745 0.610 ;
        RECT  1.945 0.275 2.055 0.610 ;
        RECT  1.255 0.510 1.945 0.610 ;
        RECT  1.145 0.275 1.255 0.610 ;
        RECT  0.455 0.510 1.145 0.610 ;
        RECT  0.345 0.275 0.455 0.610 ;
        RECT  0.150 0.510 0.345 0.610 ;
        RECT  0.050 0.510 0.150 1.305 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.4368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 0.770 3.040 0.880 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.115 -0.165 3.200 0.165 ;
        RECT  3.005 -0.165 3.115 0.445 ;
        RECT  2.625 -0.165 3.005 0.165 ;
        RECT  2.455 -0.165 2.625 0.410 ;
        RECT  2.345 -0.165 2.455 0.165 ;
        RECT  2.175 -0.165 2.345 0.410 ;
        RECT  1.825 -0.165 2.175 0.165 ;
        RECT  1.655 -0.165 1.825 0.410 ;
        RECT  1.545 -0.165 1.655 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.410 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.115 1.635 3.200 1.965 ;
        RECT  3.005 1.355 3.115 1.965 ;
        RECT  2.625 1.635 3.005 1.965 ;
        RECT  2.455 1.395 2.625 1.965 ;
        RECT  2.345 1.635 2.455 1.965 ;
        RECT  2.175 1.395 2.345 1.965 ;
        RECT  1.825 1.635 2.175 1.965 ;
        RECT  1.655 1.395 1.825 1.965 ;
        RECT  1.545 1.635 1.655 1.965 ;
        RECT  1.375 1.395 1.545 1.965 ;
        RECT  1.025 1.635 1.375 1.965 ;
        RECT  0.855 1.395 1.025 1.965 ;
        RECT  0.745 1.635 0.855 1.965 ;
        RECT  0.575 1.395 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.395 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
END GINVD8

MACRO GMUX2D1
    CLASS CORE ;
    FOREIGN GMUX2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.305 0.225 0.415 ;
        RECT  0.150 1.385 0.225 1.495 ;
        RECT  0.050 0.305 0.150 1.495 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.160 1.090 ;
        RECT  1.150 1.000 2.050 1.090 ;
        RECT  1.040 0.710 1.150 1.090 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.760 1.090 ;
        RECT  0.560 0.980 0.650 1.090 ;
        RECT  0.450 0.710 0.560 1.090 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.950 0.910 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 -0.165 2.400 0.165 ;
        RECT  1.915 -0.165 2.085 0.415 ;
        RECT  0.485 -0.165 1.915 0.165 ;
        RECT  0.315 -0.165 0.485 0.415 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 1.635 2.400 1.965 ;
        RECT  1.915 1.190 2.085 1.965 ;
        RECT  0.485 1.635 1.915 1.965 ;
        RECT  0.315 1.200 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.250 0.305 2.350 1.495 ;
        RECT  2.175 0.305 2.250 0.415 ;
        RECT  1.540 0.530 2.250 0.620 ;
        RECT  2.175 1.385 2.250 1.495 ;
        RECT  1.375 0.305 1.825 0.415 ;
        RECT  1.650 1.190 1.795 1.525 ;
        RECT  1.370 1.190 1.550 1.525 ;
        RECT  1.450 0.530 1.540 0.820 ;
        RECT  1.370 0.730 1.450 0.820 ;
        RECT  1.240 0.730 1.370 0.910 ;
        RECT  1.125 1.180 1.280 1.325 ;
        RECT  1.025 1.415 1.270 1.525 ;
        RECT  1.145 0.275 1.255 0.620 ;
        RECT  0.950 0.530 1.145 0.620 ;
        RECT  0.950 1.180 1.125 1.300 ;
        RECT  0.575 0.305 1.025 0.415 ;
        RECT  0.845 1.390 1.025 1.525 ;
        RECT  0.850 0.530 0.950 1.300 ;
        RECT  0.330 0.530 0.850 0.620 ;
        RECT  0.575 1.200 0.750 1.525 ;
        RECT  0.240 0.530 0.330 0.920 ;
        LAYER VIA1 ;
        RECT  1.650 1.250 1.750 1.350 ;
        RECT  1.410 1.190 1.510 1.290 ;
        RECT  1.110 1.415 1.210 1.515 ;
        RECT  0.650 1.290 0.750 1.390 ;
        LAYER M2 ;
        RECT  1.650 1.210 1.750 1.515 ;
        RECT  1.070 1.415 1.650 1.515 ;
        RECT  0.750 1.190 1.550 1.290 ;
        RECT  0.650 1.190 0.750 1.430 ;
    END
END GMUX2D1

MACRO GMUX2D2
    CLASS CORE ;
    FOREIGN GMUX2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.190 0.485 1.300 ;
        RECT  0.345 0.275 0.455 0.620 ;
        RECT  0.150 0.510 0.345 0.620 ;
        RECT  0.050 0.510 0.150 1.300 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.960 1.090 ;
        RECT  1.950 1.000 2.850 1.090 ;
        RECT  1.840 0.710 1.950 1.090 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.560 1.090 ;
        RECT  1.360 0.980 1.450 1.090 ;
        RECT  1.250 0.710 1.360 1.090 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.750 0.910 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.165 3.200 0.165 ;
        RECT  2.715 -0.165 2.885 0.415 ;
        RECT  1.285 -0.165 2.715 0.165 ;
        RECT  1.115 -0.165 1.285 0.415 ;
        RECT  1.025 -0.165 1.115 0.165 ;
        RECT  0.855 -0.165 1.025 0.415 ;
        RECT  0.715 -0.165 0.855 0.165 ;
        RECT  0.605 -0.165 0.715 0.445 ;
        RECT  0.225 -0.165 0.605 0.165 ;
        RECT  0.055 -0.165 0.225 0.415 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.635 3.200 1.965 ;
        RECT  2.715 1.190 2.885 1.965 ;
        RECT  1.285 1.635 2.715 1.965 ;
        RECT  1.115 1.200 1.285 1.965 ;
        RECT  0.995 1.635 1.115 1.965 ;
        RECT  0.885 1.355 0.995 1.965 ;
        RECT  0.715 1.635 0.885 1.965 ;
        RECT  0.605 1.355 0.715 1.965 ;
        RECT  0.225 1.635 0.605 1.965 ;
        RECT  0.055 1.395 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.050 0.305 3.150 1.495 ;
        RECT  2.975 0.305 3.050 0.415 ;
        RECT  2.340 0.530 3.050 0.620 ;
        RECT  2.975 1.385 3.050 1.495 ;
        RECT  2.175 0.305 2.625 0.415 ;
        RECT  2.450 1.190 2.595 1.525 ;
        RECT  2.170 1.190 2.350 1.525 ;
        RECT  2.250 0.530 2.340 0.820 ;
        RECT  2.170 0.730 2.250 0.820 ;
        RECT  2.040 0.730 2.170 0.910 ;
        RECT  1.925 1.180 2.080 1.325 ;
        RECT  1.825 1.415 2.070 1.525 ;
        RECT  1.945 0.275 2.055 0.620 ;
        RECT  1.750 0.530 1.945 0.620 ;
        RECT  1.750 1.180 1.925 1.300 ;
        RECT  1.375 0.305 1.825 0.415 ;
        RECT  1.645 1.390 1.825 1.525 ;
        RECT  1.650 0.530 1.750 1.300 ;
        RECT  0.930 0.530 1.650 0.620 ;
        RECT  1.375 1.200 1.550 1.525 ;
        RECT  1.020 0.710 1.140 1.090 ;
        RECT  0.840 0.530 0.930 0.840 ;
        RECT  0.570 0.730 0.840 0.840 ;
        RECT  0.460 0.730 0.570 0.920 ;
        RECT  0.340 0.730 0.460 0.840 ;
        RECT  0.240 0.730 0.340 0.920 ;
        LAYER VIA1 ;
        RECT  2.450 1.250 2.550 1.350 ;
        RECT  2.210 1.190 2.310 1.290 ;
        RECT  1.910 1.415 2.010 1.515 ;
        RECT  1.450 1.290 1.550 1.390 ;
        LAYER M2 ;
        RECT  2.450 1.210 2.550 1.515 ;
        RECT  1.870 1.415 2.450 1.515 ;
        RECT  1.550 1.190 2.350 1.290 ;
        RECT  1.450 1.190 1.550 1.430 ;
    END
END GMUX2D2

MACRO GMUX2ND1
    CLASS CORE ;
    FOREIGN GMUX2ND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.305 0.225 0.415 ;
        RECT  0.150 1.385 0.225 1.495 ;
        RECT  0.050 0.305 0.150 1.495 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.960 1.090 ;
        RECT  1.950 1.000 2.850 1.090 ;
        RECT  1.840 0.710 1.950 1.090 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.560 1.090 ;
        RECT  1.360 0.980 1.450 1.090 ;
        RECT  1.250 0.710 1.360 1.090 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.750 0.910 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.165 3.200 0.165 ;
        RECT  2.715 -0.165 2.885 0.415 ;
        RECT  1.285 -0.165 2.715 0.165 ;
        RECT  1.115 -0.165 1.285 0.415 ;
        RECT  0.745 -0.165 1.115 0.165 ;
        RECT  0.575 -0.165 0.745 0.415 ;
        RECT  0.000 -0.165 0.575 0.165 ;
        RECT  0.315 0.305 0.575 0.415 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.635 3.200 1.965 ;
        RECT  2.715 1.190 2.885 1.965 ;
        RECT  1.285 1.635 2.715 1.965 ;
        RECT  1.115 1.200 1.285 1.965 ;
        RECT  0.715 1.635 1.115 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.315 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.050 0.305 3.150 1.495 ;
        RECT  2.975 0.305 3.050 0.415 ;
        RECT  2.340 0.530 3.050 0.620 ;
        RECT  2.975 1.385 3.050 1.495 ;
        RECT  2.175 0.305 2.625 0.415 ;
        RECT  2.450 1.190 2.595 1.525 ;
        RECT  2.170 1.190 2.350 1.525 ;
        RECT  2.250 0.530 2.340 0.820 ;
        RECT  2.170 0.730 2.250 0.820 ;
        RECT  2.040 0.730 2.170 0.910 ;
        RECT  1.925 1.180 2.080 1.325 ;
        RECT  1.825 1.415 2.070 1.525 ;
        RECT  1.945 0.275 2.055 0.620 ;
        RECT  1.750 0.530 1.945 0.620 ;
        RECT  1.750 1.180 1.925 1.300 ;
        RECT  1.375 0.305 1.825 0.415 ;
        RECT  1.645 1.390 1.825 1.525 ;
        RECT  1.650 0.530 1.750 1.300 ;
        RECT  1.130 0.530 1.650 0.620 ;
        RECT  1.375 1.200 1.550 1.525 ;
        RECT  1.040 0.530 1.130 0.920 ;
        RECT  0.950 0.305 1.025 0.415 ;
        RECT  0.950 1.385 1.025 1.495 ;
        RECT  0.850 0.305 0.950 1.495 ;
        RECT  0.350 1.000 0.850 1.090 ;
        RECT  0.450 0.510 0.560 0.910 ;
        RECT  0.240 0.510 0.350 1.090 ;
        LAYER VIA1 ;
        RECT  2.450 1.250 2.550 1.350 ;
        RECT  2.210 1.190 2.310 1.290 ;
        RECT  1.910 1.415 2.010 1.515 ;
        RECT  1.450 1.290 1.550 1.390 ;
        LAYER M2 ;
        RECT  2.450 1.210 2.550 1.515 ;
        RECT  1.870 1.415 2.450 1.515 ;
        RECT  1.550 1.190 2.350 1.290 ;
        RECT  1.450 1.190 1.550 1.430 ;
    END
END GMUX2ND1

MACRO GMUX2ND2
    CLASS CORE ;
    FOREIGN GMUX2ND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.190 0.485 1.300 ;
        RECT  0.345 0.275 0.455 0.620 ;
        RECT  0.150 0.510 0.345 0.620 ;
        RECT  0.050 0.510 0.150 1.300 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.960 1.090 ;
        RECT  1.950 1.000 2.850 1.090 ;
        RECT  1.840 0.710 1.950 1.090 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.560 1.090 ;
        RECT  1.360 0.980 1.450 1.090 ;
        RECT  1.250 0.710 1.360 1.090 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.750 0.910 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.165 3.200 0.165 ;
        RECT  2.715 -0.165 2.885 0.415 ;
        RECT  1.285 -0.165 2.715 0.165 ;
        RECT  1.115 -0.165 1.285 0.415 ;
        RECT  0.725 -0.165 1.115 0.165 ;
        RECT  0.595 -0.165 0.725 0.465 ;
        RECT  0.225 -0.165 0.595 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.635 3.200 1.965 ;
        RECT  2.715 1.190 2.885 1.965 ;
        RECT  1.285 1.635 2.715 1.965 ;
        RECT  1.115 1.200 1.285 1.965 ;
        RECT  0.715 1.635 1.115 1.965 ;
        RECT  0.605 1.355 0.715 1.965 ;
        RECT  0.225 1.635 0.605 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.050 0.305 3.150 1.495 ;
        RECT  2.975 0.305 3.050 0.415 ;
        RECT  2.340 0.530 3.050 0.620 ;
        RECT  2.975 1.385 3.050 1.495 ;
        RECT  2.175 0.305 2.625 0.415 ;
        RECT  2.450 1.190 2.595 1.525 ;
        RECT  2.170 1.190 2.350 1.525 ;
        RECT  2.250 0.530 2.340 0.820 ;
        RECT  2.170 0.730 2.250 0.820 ;
        RECT  2.040 0.730 2.170 0.910 ;
        RECT  1.925 1.180 2.080 1.325 ;
        RECT  1.825 1.415 2.070 1.525 ;
        RECT  1.945 0.275 2.055 0.620 ;
        RECT  1.750 0.530 1.945 0.620 ;
        RECT  1.750 1.180 1.925 1.300 ;
        RECT  1.375 0.305 1.825 0.415 ;
        RECT  1.645 1.390 1.825 1.525 ;
        RECT  1.650 0.530 1.750 1.300 ;
        RECT  1.130 0.530 1.650 0.620 ;
        RECT  1.375 1.200 1.550 1.525 ;
        RECT  1.040 0.530 1.130 0.920 ;
        RECT  0.950 0.305 1.025 0.415 ;
        RECT  0.950 1.385 1.025 1.495 ;
        RECT  0.850 0.305 0.950 1.495 ;
        RECT  0.570 1.000 0.850 1.090 ;
        RECT  0.460 0.730 0.570 1.090 ;
        RECT  0.340 1.000 0.460 1.090 ;
        RECT  0.240 0.730 0.340 1.090 ;
        LAYER VIA1 ;
        RECT  2.450 1.250 2.550 1.350 ;
        RECT  2.210 1.190 2.310 1.290 ;
        RECT  1.910 1.415 2.010 1.515 ;
        RECT  1.450 1.290 1.550 1.390 ;
        LAYER M2 ;
        RECT  2.450 1.210 2.550 1.515 ;
        RECT  1.870 1.415 2.450 1.515 ;
        RECT  1.550 1.190 2.350 1.290 ;
        RECT  1.450 1.190 1.550 1.430 ;
    END
END GMUX2ND2

MACRO GND2D1
    CLASS CORE ;
    FOREIGN GND2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.275 0.750 1.300 ;
        RECT  0.605 0.275 0.650 0.560 ;
        RECT  0.315 1.190 0.650 1.300 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.690 0.560 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.690 0.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.165 0.800 0.165 ;
        RECT  0.085 -0.165 0.195 0.445 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 1.635 0.800 1.965 ;
        RECT  0.575 1.390 0.745 1.965 ;
        RECT  0.195 1.635 0.575 1.965 ;
        RECT  0.085 1.355 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.275 0.485 0.560 ;
    END
END GND2D1

MACRO GND2D2
    CLASS CORE ;
    FOREIGN GND2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.4840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.550 1.550 1.505 ;
        RECT  1.330 0.550 1.450 0.640 ;
        RECT  0.575 1.395 1.450 1.505 ;
        RECT  1.240 0.530 1.330 0.640 ;
        RECT  0.995 0.530 1.240 0.620 ;
        RECT  0.885 0.275 0.995 0.620 ;
        RECT  0.715 0.530 0.885 0.620 ;
        RECT  0.605 0.275 0.715 0.620 ;
        RECT  0.360 0.530 0.605 0.620 ;
        RECT  0.270 0.530 0.360 0.640 ;
        RECT  0.150 0.550 0.270 0.640 ;
        RECT  0.150 1.200 0.195 1.525 ;
        RECT  0.050 0.550 0.150 1.525 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.730 1.360 1.105 ;
        RECT  0.350 1.015 1.240 1.105 ;
        RECT  0.240 0.730 0.350 1.105 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.710 1.150 0.925 ;
        RECT  0.565 0.710 1.035 0.820 ;
        RECT  0.450 0.710 0.565 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 -0.165 1.600 0.165 ;
        RECT  1.415 -0.165 1.525 0.455 ;
        RECT  0.185 -0.165 1.415 0.165 ;
        RECT  0.075 -0.165 0.185 0.445 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 1.635 1.600 1.965 ;
        RECT  0.485 1.195 1.285 1.305 ;
        RECT  0.315 1.195 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.255 1.325 0.440 ;
        RECT  0.275 0.255 0.515 0.440 ;
    END
END GND2D2

MACRO GND2D3
    CLASS CORE ;
    FOREIGN GND2D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.5100 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.900 1.190 2.095 1.300 ;
        RECT  1.470 1.175 1.900 1.300 ;
        RECT  0.950 1.190 1.470 1.300 ;
        RECT  0.850 1.110 0.950 1.300 ;
        RECT  0.500 1.175 0.850 1.300 ;
        RECT  0.150 1.190 0.500 1.300 ;
        RECT  0.150 0.275 0.195 0.600 ;
        RECT  0.050 0.275 0.150 1.300 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.730 2.160 1.090 ;
        RECT  1.950 0.730 2.050 0.850 ;
        RECT  1.840 0.730 1.950 0.910 ;
        RECT  1.360 0.730 1.840 0.850 ;
        RECT  1.250 0.730 1.360 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.730 1.150 1.090 ;
        RECT  0.560 0.730 1.040 0.850 ;
        RECT  0.450 0.730 0.560 0.910 ;
        RECT  0.350 0.730 0.450 0.850 ;
        RECT  0.240 0.730 0.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 -0.165 2.400 0.165 ;
        RECT  2.205 -0.165 2.315 0.470 ;
        RECT  1.825 -0.165 2.205 0.165 ;
        RECT  1.655 -0.165 1.825 0.410 ;
        RECT  1.545 -0.165 1.655 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  0.000 -0.165 1.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 1.635 2.400 1.965 ;
        RECT  2.205 1.345 2.315 1.965 ;
        RECT  1.825 1.635 2.205 1.965 ;
        RECT  1.655 1.390 1.825 1.965 ;
        RECT  1.545 1.635 1.655 1.965 ;
        RECT  1.375 1.390 1.545 1.965 ;
        RECT  1.025 1.635 1.375 1.965 ;
        RECT  0.855 1.390 1.025 1.965 ;
        RECT  0.745 1.635 0.855 1.965 ;
        RECT  0.575 1.390 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.945 0.275 2.055 0.625 ;
        RECT  1.255 0.530 1.945 0.625 ;
        RECT  1.145 0.275 1.255 0.625 ;
        RECT  0.455 0.530 1.145 0.625 ;
        RECT  0.850 0.260 1.025 0.440 ;
        RECT  0.575 0.295 0.850 0.405 ;
        RECT  0.345 0.275 0.455 0.625 ;
        LAYER VIA1 ;
        RECT  0.850 0.300 0.950 0.400 ;
        RECT  0.850 1.150 0.950 1.250 ;
        LAYER M2 ;
        RECT  0.850 0.260 0.950 1.290 ;
    END
END GND2D3

MACRO GND2D4
    CLASS CORE ;
    FOREIGN GND2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.6800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 1.190 2.895 1.300 ;
        RECT  1.450 1.110 1.550 1.300 ;
        RECT  0.950 1.190 1.450 1.300 ;
        RECT  0.850 1.110 0.950 1.300 ;
        RECT  0.150 1.190 0.850 1.300 ;
        RECT  0.150 0.275 0.195 0.600 ;
        RECT  0.050 0.275 0.150 1.300 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.960 1.090 ;
        RECT  1.790 0.770 2.850 0.880 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.770 1.410 0.880 ;
        RECT  0.240 0.710 0.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.115 -0.165 3.200 0.165 ;
        RECT  3.005 -0.165 3.115 0.470 ;
        RECT  2.625 -0.165 3.005 0.165 ;
        RECT  2.455 -0.165 2.625 0.410 ;
        RECT  2.345 -0.165 2.455 0.165 ;
        RECT  2.175 -0.165 2.345 0.410 ;
        RECT  1.825 -0.165 2.175 0.165 ;
        RECT  1.655 -0.165 1.825 0.410 ;
        RECT  0.000 -0.165 1.655 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.115 1.635 3.200 1.965 ;
        RECT  3.005 1.345 3.115 1.965 ;
        RECT  2.625 1.635 3.005 1.965 ;
        RECT  2.455 1.390 2.625 1.965 ;
        RECT  2.345 1.635 2.455 1.965 ;
        RECT  2.175 1.390 2.345 1.965 ;
        RECT  1.825 1.635 2.175 1.965 ;
        RECT  1.655 1.390 1.825 1.965 ;
        RECT  1.545 1.635 1.655 1.965 ;
        RECT  1.375 1.390 1.545 1.965 ;
        RECT  1.025 1.635 1.375 1.965 ;
        RECT  0.855 1.390 1.025 1.965 ;
        RECT  0.745 1.635 0.855 1.965 ;
        RECT  0.575 1.390 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.145 0.275 1.255 0.660 ;
        RECT  0.750 0.550 1.145 0.660 ;
        RECT  0.850 0.260 1.025 0.440 ;
        RECT  0.575 0.295 0.850 0.405 ;
        RECT  0.640 0.520 0.750 0.660 ;
        RECT  0.455 0.520 0.640 0.620 ;
        RECT  0.345 0.275 0.455 0.620 ;
        RECT  2.745 0.275 2.855 0.620 ;
        RECT  2.560 0.520 2.745 0.620 ;
        RECT  2.450 0.520 2.560 0.660 ;
        RECT  2.055 0.550 2.450 0.660 ;
        RECT  1.945 0.275 2.055 0.660 ;
        RECT  1.255 0.550 1.945 0.660 ;
        RECT  1.345 0.260 1.565 0.460 ;
        LAYER VIA1 ;
        RECT  1.450 0.300 1.550 0.400 ;
        RECT  1.450 1.150 1.550 1.250 ;
        RECT  0.850 0.300 0.950 0.400 ;
        RECT  0.850 1.150 0.950 1.250 ;
        LAYER M2 ;
        RECT  1.450 0.260 1.550 1.290 ;
        RECT  0.850 0.260 0.950 1.290 ;
    END
END GND2D4

MACRO GND3D1
    CLASS CORE ;
    FOREIGN GND3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2580 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.885 1.190 0.995 1.525 ;
        RECT  0.150 1.190 0.885 1.300 ;
        RECT  0.150 0.275 0.195 0.550 ;
        RECT  0.050 0.275 0.150 1.300 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.690 0.350 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.570 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.690 1.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 -0.165 1.600 0.165 ;
        RECT  1.405 -0.165 1.515 0.445 ;
        RECT  1.255 -0.165 1.405 0.165 ;
        RECT  1.145 -0.165 1.255 0.445 ;
        RECT  0.000 -0.165 1.145 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.200 1.515 1.965 ;
        RECT  1.115 1.200 1.405 1.310 ;
        RECT  0.360 1.635 1.405 1.965 ;
        RECT  0.360 1.390 0.745 1.500 ;
        RECT  0.240 1.390 0.360 1.965 ;
        RECT  0.055 1.390 0.240 1.500 ;
        RECT  0.000 1.635 0.240 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.740 1.500 0.930 ;
        RECT  0.575 0.305 1.025 0.415 ;
        RECT  0.315 0.275 0.485 0.550 ;
    END
END GND3D1

MACRO GND3D2
    CLASS CORE ;
    FOREIGN GND3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.4440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.275 2.350 1.300 ;
        RECT  2.205 0.275 2.250 0.600 ;
        RECT  0.150 1.195 2.250 1.300 ;
        RECT  0.150 0.275 0.195 0.600 ;
        RECT  0.050 0.275 0.150 1.300 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.710 1.370 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.730 1.950 0.920 ;
        RECT  1.650 0.510 1.750 0.920 ;
        RECT  0.750 0.510 1.650 0.610 ;
        RECT  0.650 0.510 0.750 0.920 ;
        RECT  0.450 0.730 0.650 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.710 2.160 1.105 ;
        RECT  0.350 1.015 2.040 1.105 ;
        RECT  0.240 0.710 0.350 1.105 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 -0.165 2.400 0.165 ;
        RECT  1.115 -0.165 1.285 0.415 ;
        RECT  0.000 -0.165 1.115 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.635 2.400 1.965 ;
        RECT  2.175 1.390 2.345 1.965 ;
        RECT  1.825 1.635 2.175 1.965 ;
        RECT  1.655 1.390 1.825 1.965 ;
        RECT  1.545 1.635 1.655 1.965 ;
        RECT  1.375 1.390 1.545 1.965 ;
        RECT  1.025 1.635 1.375 1.965 ;
        RECT  0.855 1.390 1.025 1.965 ;
        RECT  0.745 1.635 0.855 1.965 ;
        RECT  0.575 1.390 0.745 1.965 ;
        RECT  0.225 1.635 0.575 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.275 2.075 0.600 ;
        RECT  1.375 0.305 1.825 0.415 ;
        RECT  0.575 0.305 1.025 0.415 ;
        RECT  0.325 0.275 0.475 0.600 ;
    END
END GND3D2

MACRO GNR2D1
    CLASS CORE ;
    FOREIGN GNR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1660 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.500 0.750 1.525 ;
        RECT  0.455 0.500 0.650 0.600 ;
        RECT  0.600 1.210 0.650 1.525 ;
        RECT  0.345 0.275 0.455 0.600 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.690 0.560 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.690 0.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 0.800 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.195 -0.165 0.575 0.165 ;
        RECT  0.085 -0.165 0.195 0.445 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.635 0.800 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 1.200 0.490 1.350 ;
        RECT  0.070 1.200 0.315 1.300 ;
    END
END GNR2D1

MACRO GNR2D2
    CLASS CORE ;
    FOREIGN GNR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.525 ;
        RECT  1.255 0.510 1.450 0.620 ;
        RECT  1.405 1.200 1.450 1.525 ;
        RECT  1.145 0.275 1.255 0.620 ;
        RECT  0.455 0.530 1.145 0.620 ;
        RECT  0.345 0.275 0.455 0.620 ;
        RECT  0.150 0.510 0.345 0.620 ;
        RECT  0.150 1.200 0.195 1.525 ;
        RECT  0.050 0.510 0.150 1.525 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.710 1.360 1.105 ;
        RECT  0.360 1.015 1.240 1.105 ;
        RECT  0.240 0.710 0.360 1.105 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.710 1.150 0.925 ;
        RECT  0.565 0.710 1.035 0.820 ;
        RECT  0.450 0.710 0.565 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.420 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.420 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.420 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.420 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.635 1.600 1.965 ;
        RECT  0.760 1.395 1.025 1.505 ;
        RECT  0.640 1.395 0.760 1.965 ;
        RECT  0.575 1.395 0.640 1.505 ;
        RECT  0.000 1.635 0.640 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.115 1.195 1.285 1.505 ;
        RECT  0.315 1.195 0.485 1.505 ;
    END
END GNR2D2

MACRO GNR3D1
    CLASS CORE ;
    FOREIGN GNR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.885 0.275 0.995 0.600 ;
        RECT  0.455 0.500 0.885 0.600 ;
        RECT  0.345 0.275 0.455 0.600 ;
        RECT  0.150 0.500 0.345 0.600 ;
        RECT  0.150 1.355 0.225 1.525 ;
        RECT  0.050 0.500 0.150 1.525 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.690 1.150 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.690 0.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.415 ;
        RECT  0.745 -0.165 1.375 0.165 ;
        RECT  1.115 0.305 1.375 0.415 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.210 1.515 1.965 ;
        RECT  1.115 1.210 1.405 1.320 ;
        RECT  0.000 1.635 1.405 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.610 1.460 0.910 ;
        RECT  0.575 1.385 1.025 1.495 ;
        RECT  0.315 1.200 0.485 1.515 ;
    END
END GNR3D1

MACRO GNR3D2
    CLASS CORE ;
    FOREIGN GNR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.4100 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 0.275 2.055 0.600 ;
        RECT  1.255 0.500 1.945 0.600 ;
        RECT  1.145 0.275 1.255 0.600 ;
        RECT  0.455 0.500 1.145 0.600 ;
        RECT  0.150 1.390 0.745 1.500 ;
        RECT  0.345 0.275 0.455 0.600 ;
        RECT  0.150 0.500 0.345 0.600 ;
        RECT  0.050 0.500 0.150 1.500 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.690 2.160 1.090 ;
        RECT  1.950 0.980 2.050 1.090 ;
        RECT  1.840 0.690 1.950 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.690 1.360 1.090 ;
        RECT  1.150 0.980 1.250 1.090 ;
        RECT  1.040 0.690 1.150 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.690 0.560 1.090 ;
        RECT  0.350 0.980 0.450 1.090 ;
        RECT  0.240 0.690 0.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 -0.165 2.400 0.165 ;
        RECT  2.175 -0.165 2.345 0.410 ;
        RECT  1.825 -0.165 2.175 0.165 ;
        RECT  1.655 -0.165 1.825 0.410 ;
        RECT  1.545 -0.165 1.655 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.410 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.225 -0.165 0.575 0.165 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.635 2.400 1.965 ;
        RECT  2.175 1.390 2.345 1.965 ;
        RECT  1.825 1.635 2.175 1.965 ;
        RECT  1.655 1.390 1.825 1.965 ;
        RECT  0.000 1.635 1.655 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.105 1.200 2.095 1.300 ;
        RECT  0.955 1.390 1.545 1.500 ;
        RECT  0.855 1.200 0.955 1.500 ;
        RECT  0.315 1.200 0.855 1.300 ;
    END
END GNR3D2

MACRO GOAI21D1
    CLASS CORE ;
    FOREIGN GOAI21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.395 1.025 1.525 ;
        RECT  0.750 1.305 0.950 1.525 ;
        RECT  0.650 0.275 0.750 1.525 ;
        RECT  0.615 0.275 0.650 0.610 ;
        RECT  0.575 1.395 0.650 1.525 ;
        RECT  0.185 0.520 0.615 0.610 ;
        RECT  0.150 0.275 0.185 0.610 ;
        RECT  0.050 0.275 0.150 1.090 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.690 1.150 1.095 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.350 1.095 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.560 1.095 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.415 ;
        RECT  0.000 -0.165 1.375 0.165 ;
        RECT  1.115 0.305 1.375 0.415 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.210 1.515 1.965 ;
        RECT  1.115 1.210 1.405 1.320 ;
        RECT  0.225 1.635 1.405 1.965 ;
        RECT  0.055 1.375 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.610 1.460 0.910 ;
        RECT  0.850 0.275 1.005 0.580 ;
        RECT  0.275 0.255 0.525 0.430 ;
        RECT  0.315 1.205 0.485 1.525 ;
        LAYER VIA1 ;
        RECT  0.850 0.350 0.950 0.450 ;
        RECT  0.350 0.310 0.450 0.410 ;
        LAYER M2 ;
        RECT  0.850 0.310 0.950 0.490 ;
        RECT  0.310 0.310 0.850 0.410 ;
    END
END GOAI21D1

MACRO GOAI21D2
    CLASS CORE ;
    FOREIGN GOAI21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.5440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.275 2.350 1.525 ;
        RECT  2.210 0.275 2.250 0.615 ;
        RECT  2.195 1.300 2.250 1.525 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.560 1.095 ;
        RECT  0.350 0.985 0.450 1.095 ;
        RECT  0.240 0.710 0.350 1.095 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.710 1.950 0.910 ;
        RECT  1.360 0.800 1.840 0.910 ;
        RECT  1.250 0.710 1.360 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.160 1.115 ;
        RECT  1.150 1.020 2.050 1.115 ;
        RECT  1.040 0.710 1.150 1.115 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 2.400 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.205 -0.165 0.575 0.165 ;
        RECT  0.075 -0.165 0.205 0.445 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 1.635 2.400 1.965 ;
        RECT  1.685 1.345 1.795 1.965 ;
        RECT  1.515 1.635 1.685 1.965 ;
        RECT  1.405 1.345 1.515 1.965 ;
        RECT  0.745 1.635 1.405 1.965 ;
        RECT  0.575 1.390 0.745 1.965 ;
        RECT  0.205 1.635 0.575 1.965 ;
        RECT  0.075 1.355 0.205 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.090 0.275 2.095 0.375 ;
        RECT  1.910 0.275 2.090 0.580 ;
        RECT  1.915 1.210 2.085 1.525 ;
        RECT  1.655 0.275 1.785 0.580 ;
        RECT  1.545 0.475 1.655 0.580 ;
        RECT  1.415 0.275 1.545 0.580 ;
        RECT  1.290 0.275 1.295 0.375 ;
        RECT  1.110 0.275 1.290 0.580 ;
        RECT  1.115 1.210 1.285 1.525 ;
        RECT  0.875 1.210 1.005 1.525 ;
        RECT  0.855 0.275 0.985 0.600 ;
        RECT  0.750 0.500 0.855 0.600 ;
        RECT  0.650 0.500 0.750 1.300 ;
        RECT  0.305 1.210 0.650 1.300 ;
        RECT  0.305 0.275 0.485 0.580 ;
        RECT  0.750 1.210 0.875 1.300 ;
        LAYER VIA1 ;
        RECT  2.210 0.475 2.310 0.575 ;
        RECT  1.955 0.275 2.055 0.375 ;
        RECT  1.550 0.475 1.650 0.575 ;
        RECT  1.155 0.275 1.255 0.375 ;
        RECT  0.650 0.540 0.750 0.640 ;
        RECT  0.345 0.275 0.445 0.375 ;
        LAYER M2 ;
        RECT  2.250 0.475 2.350 0.690 ;
        RECT  0.750 0.475 2.250 0.575 ;
        RECT  0.305 0.275 2.095 0.375 ;
        RECT  0.650 0.475 0.750 0.680 ;
    END
END GOAI21D2

MACRO GOR2D1
    CLASS CORE ;
    FOREIGN GOR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 0.495 1.550 1.525 ;
        RECT  1.450 0.275 1.515 1.525 ;
        RECT  1.405 0.275 1.450 0.585 ;
        RECT  1.405 1.240 1.450 1.525 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.690 0.350 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.690 0.560 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.025 -0.165 1.600 0.165 ;
        RECT  1.025 0.305 1.285 0.415 ;
        RECT  0.855 -0.165 1.025 0.415 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.195 -0.165 0.575 0.165 ;
        RECT  0.085 -0.165 0.195 0.445 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.995 1.635 1.600 1.965 ;
        RECT  0.995 1.210 1.285 1.320 ;
        RECT  0.885 1.210 0.995 1.965 ;
        RECT  0.225 1.635 0.885 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.730 1.360 1.110 ;
        RECT  0.750 1.000 1.250 1.110 ;
        RECT  0.940 0.610 1.140 0.910 ;
        RECT  0.720 0.500 0.750 1.330 ;
        RECT  0.650 0.500 0.720 1.525 ;
        RECT  0.455 0.500 0.650 0.600 ;
        RECT  0.600 1.210 0.650 1.525 ;
        RECT  0.315 1.200 0.490 1.350 ;
        RECT  0.345 0.275 0.455 0.600 ;
        RECT  0.070 1.200 0.315 1.300 ;
    END
END GOR2D1

MACRO GOR2D2
    CLASS CORE ;
    FOREIGN GOR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.300 ;
        RECT  1.255 0.510 1.450 0.630 ;
        RECT  1.105 1.190 1.450 1.300 ;
        RECT  1.145 0.275 1.255 0.630 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.690 0.350 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.690 0.560 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.165 1.600 0.165 ;
        RECT  1.375 -0.165 1.545 0.410 ;
        RECT  1.025 -0.165 1.375 0.165 ;
        RECT  0.855 -0.165 1.025 0.415 ;
        RECT  0.745 -0.165 0.855 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.195 -0.165 0.575 0.165 ;
        RECT  0.085 -0.165 0.195 0.445 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.635 1.600 1.965 ;
        RECT  1.375 1.390 1.545 1.965 ;
        RECT  0.995 1.635 1.375 1.965 ;
        RECT  0.885 1.355 0.995 1.965 ;
        RECT  0.225 1.635 0.885 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.740 1.360 1.080 ;
        RECT  1.140 0.970 1.250 1.080 ;
        RECT  1.030 0.740 1.140 1.080 ;
        RECT  0.750 0.970 1.030 1.080 ;
        RECT  0.720 0.500 0.750 1.330 ;
        RECT  0.650 0.500 0.720 1.525 ;
        RECT  0.455 0.500 0.650 0.600 ;
        RECT  0.600 1.210 0.650 1.525 ;
        RECT  0.315 1.200 0.490 1.350 ;
        RECT  0.345 0.275 0.455 0.600 ;
        RECT  0.070 1.200 0.315 1.300 ;
    END
END GOR2D2

MACRO GSDFCNQD1
    CLASS CORE ;
    FOREIGN GSDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN SI
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.710 0.350 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.780 1.170 0.890 ;
        RECT  0.440 0.710 0.560 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.305 7.150 1.495 ;
        RECT  6.975 0.305 7.050 0.415 ;
        RECT  6.975 1.385 7.050 1.495 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.510 1.955 0.910 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.540 4.560 0.910 ;
        RECT  3.150 0.540 4.450 0.630 ;
        RECT  3.040 0.510 3.150 0.910 ;
        RECT  2.850 0.710 3.040 0.910 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  3.950 1.010 5.945 1.110 ;
        RECT  3.850 0.730 3.950 1.110 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.865 -0.165 7.200 0.165 ;
        RECT  6.735 -0.165 6.865 0.495 ;
        RECT  5.790 -0.165 6.735 0.165 ;
        RECT  5.680 -0.165 5.790 0.445 ;
        RECT  4.465 -0.165 5.680 0.165 ;
        RECT  4.335 -0.165 4.465 0.445 ;
        RECT  3.930 -0.165 4.335 0.165 ;
        RECT  3.815 -0.165 3.930 0.450 ;
        RECT  2.085 -0.165 3.815 0.165 ;
        RECT  1.915 -0.165 2.085 0.415 ;
        RECT  0.455 -0.165 1.915 0.165 ;
        RECT  0.345 -0.165 0.455 0.465 ;
        RECT  0.000 -0.165 0.345 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.870 1.635 7.200 1.965 ;
        RECT  6.735 1.150 6.870 1.965 ;
        RECT  6.085 1.635 6.735 1.965 ;
        RECT  5.915 1.210 6.085 1.965 ;
        RECT  4.485 1.635 5.915 1.965 ;
        RECT  4.315 1.210 4.485 1.965 ;
        RECT  3.685 1.635 4.315 1.965 ;
        RECT  3.515 1.210 3.685 1.965 ;
        RECT  2.085 1.635 3.515 1.965 ;
        RECT  1.915 1.210 2.085 1.965 ;
        RECT  0.485 1.635 1.915 1.965 ;
        RECT  0.315 1.210 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.360 0.740 6.960 0.910 ;
        RECT  6.450 1.210 6.630 1.525 ;
        RECT  6.450 0.255 6.615 0.630 ;
        RECT  6.270 0.295 6.360 1.525 ;
        RECT  6.175 0.295 6.270 0.420 ;
        RECT  6.180 1.210 6.270 1.525 ;
        RECT  6.030 0.600 6.170 1.110 ;
        RECT  5.905 0.255 6.085 0.490 ;
        RECT  5.745 1.010 6.030 1.110 ;
        RECT  5.635 0.740 5.930 0.910 ;
        RECT  5.635 1.215 5.815 1.525 ;
        RECT  5.545 0.540 5.635 1.110 ;
        RECT  5.345 0.255 5.590 0.450 ;
        RECT  5.255 0.540 5.545 0.630 ;
        RECT  5.255 1.010 5.545 1.110 ;
        RECT  5.380 1.210 5.525 1.525 ;
        RECT  5.220 0.720 5.440 0.920 ;
        RECT  5.145 0.275 5.255 0.630 ;
        RECT  5.145 1.010 5.255 1.360 ;
        RECT  4.750 0.740 5.130 0.910 ;
        RECT  4.850 0.255 5.035 0.650 ;
        RECT  4.850 1.210 5.020 1.510 ;
        RECT  4.650 0.300 4.750 1.505 ;
        RECT  4.575 0.300 4.650 0.425 ;
        RECT  4.575 1.380 4.650 1.505 ;
        RECT  4.230 0.730 4.340 1.110 ;
        RECT  4.020 0.255 4.245 0.450 ;
        RECT  2.855 1.010 4.230 1.110 ;
        RECT  4.050 1.210 4.220 1.510 ;
        RECT  3.775 1.210 3.955 1.510 ;
        RECT  3.650 0.730 3.950 0.910 ;
        RECT  3.505 0.255 3.725 0.450 ;
        RECT  3.315 0.740 3.550 0.920 ;
        RECT  3.245 1.210 3.425 1.510 ;
        RECT  3.250 0.275 3.395 0.445 ;
        RECT  2.955 0.275 3.250 0.405 ;
        RECT  2.965 1.210 3.145 1.510 ;
        RECT  2.745 0.255 2.865 0.610 ;
        RECT  2.745 1.010 2.855 1.350 ;
        RECT  2.675 1.010 2.745 1.110 ;
        RECT  2.555 0.740 2.740 0.910 ;
        RECT  2.410 0.255 2.655 0.460 ;
        RECT  2.450 1.220 2.630 1.510 ;
        RECT  2.465 0.550 2.555 1.110 ;
        RECT  2.320 0.550 2.465 0.640 ;
        RECT  2.310 1.020 2.465 1.110 ;
        RECT  2.045 0.730 2.355 0.930 ;
        RECT  2.210 0.275 2.320 0.640 ;
        RECT  2.205 1.020 2.310 1.525 ;
        RECT  1.745 0.305 1.825 0.415 ;
        RECT  1.745 1.385 1.825 1.495 ;
        RECT  1.650 0.305 1.745 1.495 ;
        RECT  1.375 0.305 1.650 0.415 ;
        RECT  1.565 1.010 1.650 1.110 ;
        RECT  1.380 1.210 1.560 1.525 ;
        RECT  1.270 0.600 1.360 1.070 ;
        RECT  1.105 1.210 1.285 1.525 ;
        RECT  1.105 0.255 1.275 0.510 ;
        RECT  0.745 0.600 1.270 0.690 ;
        RECT  0.750 0.980 1.270 1.070 ;
        RECT  0.835 0.255 1.015 0.510 ;
        RECT  0.850 1.160 0.990 1.525 ;
        RECT  0.650 0.980 0.750 1.525 ;
        RECT  0.655 0.275 0.745 0.690 ;
        RECT  0.600 0.275 0.655 0.465 ;
        RECT  0.610 1.310 0.650 1.525 ;
        RECT  0.075 0.255 0.255 0.570 ;
        RECT  0.045 1.210 0.225 1.525 ;
        LAYER VIA1 ;
        RECT  6.490 1.210 6.590 1.310 ;
        RECT  6.450 0.390 6.550 0.490 ;
        RECT  6.220 1.410 6.320 1.510 ;
        RECT  5.785 1.010 5.885 1.110 ;
        RECT  5.675 1.410 5.775 1.510 ;
        RECT  5.420 0.340 5.520 0.440 ;
        RECT  5.415 1.250 5.515 1.350 ;
        RECT  5.295 0.750 5.395 0.850 ;
        RECT  4.890 0.550 4.990 0.650 ;
        RECT  4.850 1.250 4.950 1.350 ;
        RECT  4.450 0.710 4.550 0.810 ;
        RECT  4.080 1.250 4.180 1.350 ;
        RECT  4.070 0.340 4.170 0.440 ;
        RECT  3.850 0.770 3.950 0.870 ;
        RECT  3.815 1.410 3.915 1.510 ;
        RECT  3.450 0.780 3.550 0.880 ;
        RECT  3.285 1.410 3.385 1.510 ;
        RECT  3.005 1.210 3.105 1.310 ;
        RECT  2.850 0.770 2.950 0.870 ;
        RECT  2.755 0.470 2.855 0.570 ;
        RECT  2.715 1.010 2.815 1.110 ;
        RECT  2.490 1.410 2.590 1.510 ;
        RECT  2.480 0.310 2.580 0.410 ;
        RECT  2.255 0.770 2.355 0.870 ;
        RECT  1.605 1.010 1.705 1.110 ;
        RECT  1.420 1.410 1.520 1.510 ;
        RECT  1.155 0.310 1.255 0.410 ;
        RECT  1.145 1.210 1.245 1.310 ;
        RECT  0.875 0.310 0.975 0.410 ;
        RECT  0.850 1.200 0.950 1.300 ;
        RECT  0.115 0.310 0.215 0.410 ;
        RECT  0.085 1.390 0.185 1.490 ;
        LAYER M2 ;
        RECT  6.550 1.210 6.630 1.310 ;
        RECT  6.450 0.350 6.550 1.310 ;
        RECT  5.850 0.350 6.450 0.450 ;
        RECT  5.515 1.210 6.450 1.310 ;
        RECT  5.635 1.410 6.360 1.510 ;
        RECT  5.750 0.350 5.850 0.650 ;
        RECT  4.850 0.550 5.750 0.650 ;
        RECT  3.550 0.340 5.560 0.440 ;
        RECT  5.415 1.210 5.515 1.390 ;
        RECT  4.550 0.750 5.435 0.850 ;
        RECT  4.850 1.210 4.950 1.390 ;
        RECT  4.180 1.210 4.850 1.310 ;
        RECT  4.450 0.670 4.550 0.850 ;
        RECT  4.080 1.210 4.180 1.390 ;
        RECT  3.550 1.210 4.080 1.310 ;
        RECT  2.450 1.410 3.955 1.510 ;
        RECT  3.450 0.340 3.550 1.310 ;
        RECT  1.105 1.210 3.145 1.310 ;
        RECT  2.850 0.730 2.950 0.910 ;
        RECT  2.755 0.430 2.855 0.610 ;
        RECT  2.150 1.010 2.855 1.110 ;
        RECT  2.355 0.810 2.850 0.910 ;
        RECT  2.150 0.510 2.755 0.610 ;
        RECT  1.115 0.310 2.620 0.410 ;
        RECT  2.255 0.730 2.355 0.910 ;
        RECT  2.050 0.510 2.150 1.110 ;
        RECT  0.950 1.010 1.745 1.110 ;
        RECT  1.380 1.410 1.560 1.540 ;
        RECT  0.205 1.440 1.380 1.540 ;
        RECT  0.075 0.310 1.015 0.410 ;
        RECT  0.850 1.010 0.950 1.340 ;
        RECT  0.065 1.340 0.205 1.540 ;
    END
END GSDFCNQD1

MACRO GTIEH
    CLASS CORE ;
    FOREIGN GTIEH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.0880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.200 0.195 1.525 ;
        RECT  0.050 0.710 0.150 1.525 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 0.800 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.485 -0.165 0.575 0.165 ;
        RECT  0.315 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.315 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.450 0.710 0.570 1.090 ;
        RECT  0.240 0.510 0.360 0.910 ;
        RECT  0.195 0.510 0.240 0.600 ;
        RECT  0.085 0.265 0.195 0.600 ;
    END
END GTIEH

MACRO GTIEL
    CLASS CORE ;
    FOREIGN GTIEL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.265 0.195 0.455 ;
        RECT  0.050 0.265 0.150 0.910 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 0.800 0.165 ;
        RECT  0.575 -0.165 0.745 0.410 ;
        RECT  0.485 -0.165 0.575 0.165 ;
        RECT  0.315 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.200 0.715 1.965 ;
        RECT  0.315 1.200 0.605 1.310 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.450 0.710 0.570 1.090 ;
        RECT  0.240 0.710 0.360 1.110 ;
        RECT  0.195 1.020 0.240 1.110 ;
        RECT  0.085 1.020 0.195 1.525 ;
    END
END GTIEL

MACRO GXNR2D1
    CLASS CORE ;
    FOREIGN GXNR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.305 0.225 0.415 ;
        RECT  0.150 1.385 0.225 1.495 ;
        RECT  0.050 0.305 0.150 1.495 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.560 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.160 1.090 ;
        RECT  1.150 1.000 2.050 1.090 ;
        RECT  1.040 0.710 1.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 -0.165 2.400 0.165 ;
        RECT  1.915 -0.165 2.085 0.415 ;
        RECT  0.485 -0.165 1.915 0.165 ;
        RECT  0.315 -0.165 0.485 0.415 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 1.635 2.400 1.965 ;
        RECT  1.915 1.190 2.085 1.965 ;
        RECT  0.485 1.635 1.915 1.965 ;
        RECT  0.315 1.200 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.250 0.305 2.350 1.495 ;
        RECT  2.175 0.305 2.250 0.415 ;
        RECT  1.540 0.530 2.250 0.620 ;
        RECT  2.175 1.385 2.250 1.495 ;
        RECT  1.650 0.710 1.950 0.910 ;
        RECT  1.375 0.305 1.825 0.415 ;
        RECT  1.640 1.190 1.820 1.525 ;
        RECT  1.370 1.190 1.550 1.525 ;
        RECT  1.450 0.530 1.540 0.820 ;
        RECT  1.370 0.730 1.450 0.820 ;
        RECT  1.240 0.730 1.370 0.910 ;
        RECT  1.125 1.180 1.280 1.325 ;
        RECT  1.025 1.415 1.270 1.525 ;
        RECT  1.145 0.275 1.255 0.620 ;
        RECT  0.950 0.530 1.145 0.620 ;
        RECT  0.950 1.180 1.125 1.300 ;
        RECT  0.750 0.305 1.025 0.415 ;
        RECT  0.845 1.390 1.025 1.525 ;
        RECT  0.850 0.530 0.950 1.300 ;
        RECT  0.650 0.305 0.750 0.900 ;
        RECT  0.575 1.200 0.750 1.525 ;
        RECT  0.575 0.305 0.650 0.415 ;
        RECT  0.240 0.730 0.330 1.100 ;
        RECT  0.330 1.010 0.850 1.100 ;
        LAYER VIA1 ;
        RECT  1.680 1.415 1.780 1.515 ;
        RECT  1.650 0.750 1.750 0.850 ;
        RECT  1.410 1.190 1.510 1.290 ;
        RECT  1.110 1.415 1.210 1.515 ;
        RECT  0.650 0.750 0.750 0.850 ;
        RECT  0.650 1.290 0.750 1.390 ;
        LAYER M2 ;
        RECT  1.070 1.415 1.820 1.515 ;
        RECT  1.650 0.710 1.750 1.290 ;
        RECT  0.750 1.190 1.650 1.290 ;
        RECT  0.650 0.710 0.750 1.430 ;
    END
END GXNR2D1

MACRO GXNR2D2
    CLASS CORE ;
    FOREIGN GXNR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.190 0.485 1.300 ;
        RECT  0.345 0.275 0.455 0.620 ;
        RECT  0.150 0.510 0.345 0.620 ;
        RECT  0.050 0.510 0.150 1.300 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.360 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.960 1.090 ;
        RECT  1.950 1.000 2.850 1.090 ;
        RECT  1.840 0.710 1.950 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.165 3.200 0.165 ;
        RECT  2.715 -0.165 2.885 0.415 ;
        RECT  1.025 -0.165 2.715 0.165 ;
        RECT  1.025 0.305 1.285 0.415 ;
        RECT  0.855 -0.165 1.025 0.415 ;
        RECT  0.225 -0.165 0.855 0.165 ;
        RECT  0.575 0.305 0.855 0.415 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.635 3.200 1.965 ;
        RECT  2.715 1.190 2.885 1.965 ;
        RECT  0.995 1.635 2.715 1.965 ;
        RECT  0.995 1.200 1.285 1.310 ;
        RECT  0.885 1.200 0.995 1.965 ;
        RECT  0.715 1.635 0.885 1.965 ;
        RECT  0.605 1.355 0.715 1.965 ;
        RECT  0.225 1.635 0.605 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.050 0.305 3.150 1.495 ;
        RECT  2.975 0.305 3.050 0.415 ;
        RECT  2.340 0.530 3.050 0.620 ;
        RECT  2.975 1.385 3.050 1.495 ;
        RECT  2.450 0.710 2.750 0.910 ;
        RECT  2.175 0.305 2.625 0.415 ;
        RECT  2.440 1.190 2.620 1.525 ;
        RECT  2.170 1.190 2.350 1.525 ;
        RECT  2.250 0.530 2.340 0.820 ;
        RECT  2.170 0.730 2.250 0.820 ;
        RECT  2.040 0.730 2.170 0.910 ;
        RECT  1.925 1.180 2.080 1.325 ;
        RECT  1.825 1.415 2.070 1.525 ;
        RECT  1.945 0.275 2.055 0.620 ;
        RECT  1.750 0.530 1.945 0.620 ;
        RECT  1.750 1.180 1.925 1.300 ;
        RECT  1.550 0.305 1.825 0.415 ;
        RECT  1.645 1.390 1.825 1.525 ;
        RECT  1.650 0.530 1.750 1.300 ;
        RECT  0.570 1.010 1.650 1.100 ;
        RECT  1.450 0.305 1.550 0.900 ;
        RECT  1.375 1.200 1.550 1.525 ;
        RECT  1.375 0.305 1.450 0.415 ;
        RECT  1.030 0.510 1.140 0.910 ;
        RECT  0.460 0.730 0.570 1.100 ;
        RECT  0.340 1.010 0.460 1.100 ;
        RECT  0.240 0.730 0.340 1.100 ;
        LAYER VIA1 ;
        RECT  2.480 1.415 2.580 1.515 ;
        RECT  2.450 0.750 2.550 0.850 ;
        RECT  2.210 1.190 2.310 1.290 ;
        RECT  1.910 1.415 2.010 1.515 ;
        RECT  1.450 0.750 1.550 0.850 ;
        RECT  1.450 1.290 1.550 1.390 ;
        LAYER M2 ;
        RECT  1.870 1.415 2.620 1.515 ;
        RECT  2.450 0.710 2.550 1.290 ;
        RECT  1.550 1.190 2.450 1.290 ;
        RECT  1.450 0.710 1.550 1.430 ;
    END
END GXNR2D2

MACRO GXOR2D1
    CLASS CORE ;
    FOREIGN GXOR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.305 0.225 0.415 ;
        RECT  0.150 1.385 0.225 1.495 ;
        RECT  0.050 0.305 0.150 1.495 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.560 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.510 2.160 0.910 ;
        RECT  1.550 0.510 2.050 0.620 ;
        RECT  1.450 0.510 1.550 0.910 ;
        RECT  1.250 0.730 1.450 0.910 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 -0.165 2.400 0.165 ;
        RECT  1.915 -0.165 2.085 0.415 ;
        RECT  0.485 -0.165 1.915 0.165 ;
        RECT  0.315 -0.165 0.485 0.415 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 1.635 2.400 1.965 ;
        RECT  1.915 1.190 2.085 1.965 ;
        RECT  0.485 1.635 1.915 1.965 ;
        RECT  0.315 1.200 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.250 0.305 2.350 1.495 ;
        RECT  2.175 0.305 2.250 0.415 ;
        RECT  1.150 1.000 2.250 1.090 ;
        RECT  2.175 1.385 2.250 1.495 ;
        RECT  1.650 0.710 1.950 0.910 ;
        RECT  1.375 0.305 1.825 0.415 ;
        RECT  1.640 1.190 1.820 1.525 ;
        RECT  1.370 1.190 1.550 1.525 ;
        RECT  1.125 1.180 1.280 1.325 ;
        RECT  1.025 1.415 1.270 1.525 ;
        RECT  1.145 0.275 1.255 0.625 ;
        RECT  1.040 0.715 1.150 1.090 ;
        RECT  0.950 0.525 1.145 0.625 ;
        RECT  0.950 1.180 1.125 1.300 ;
        RECT  0.750 0.305 1.025 0.415 ;
        RECT  0.850 0.525 0.950 1.300 ;
        RECT  0.330 1.010 0.850 1.100 ;
        RECT  0.650 0.305 0.750 0.900 ;
        RECT  0.575 1.200 0.750 1.525 ;
        RECT  0.575 0.305 0.650 0.415 ;
        RECT  0.240 0.730 0.330 1.100 ;
        RECT  0.845 1.390 1.025 1.525 ;
        LAYER VIA1 ;
        RECT  1.680 1.415 1.780 1.515 ;
        RECT  1.650 0.750 1.750 0.850 ;
        RECT  1.410 1.190 1.510 1.290 ;
        RECT  1.110 1.415 1.210 1.515 ;
        RECT  0.650 0.750 0.750 0.850 ;
        RECT  0.650 1.290 0.750 1.390 ;
        LAYER M2 ;
        RECT  1.070 1.415 1.820 1.515 ;
        RECT  1.650 0.710 1.750 1.290 ;
        RECT  0.750 1.190 1.650 1.290 ;
        RECT  0.650 0.710 0.750 1.430 ;
    END
END GXOR2D1

MACRO GXOR2D2
    CLASS CORE ;
    FOREIGN GXOR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.190 0.485 1.300 ;
        RECT  0.345 0.275 0.455 0.620 ;
        RECT  0.150 0.510 0.345 0.620 ;
        RECT  0.050 0.510 0.150 1.300 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.360 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.510 2.960 0.910 ;
        RECT  2.350 0.510 2.850 0.620 ;
        RECT  2.250 0.510 2.350 0.910 ;
        RECT  2.050 0.730 2.250 0.910 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.165 3.200 0.165 ;
        RECT  2.715 -0.165 2.885 0.415 ;
        RECT  1.025 -0.165 2.715 0.165 ;
        RECT  1.025 0.305 1.285 0.415 ;
        RECT  0.855 -0.165 1.025 0.415 ;
        RECT  0.225 -0.165 0.855 0.165 ;
        RECT  0.575 0.305 0.855 0.415 ;
        RECT  0.055 -0.165 0.225 0.410 ;
        RECT  0.000 -0.165 0.055 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.635 3.200 1.965 ;
        RECT  2.715 1.190 2.885 1.965 ;
        RECT  0.995 1.635 2.715 1.965 ;
        RECT  0.995 1.200 1.285 1.310 ;
        RECT  0.885 1.200 0.995 1.965 ;
        RECT  0.715 1.635 0.885 1.965 ;
        RECT  0.605 1.355 0.715 1.965 ;
        RECT  0.225 1.635 0.605 1.965 ;
        RECT  0.055 1.390 0.225 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.050 0.305 3.150 1.495 ;
        RECT  2.975 0.305 3.050 0.415 ;
        RECT  1.950 1.000 3.050 1.090 ;
        RECT  2.975 1.385 3.050 1.495 ;
        RECT  2.450 0.710 2.750 0.910 ;
        RECT  2.175 0.305 2.625 0.415 ;
        RECT  2.440 1.190 2.620 1.525 ;
        RECT  2.170 1.190 2.350 1.525 ;
        RECT  1.925 1.180 2.080 1.325 ;
        RECT  1.825 1.415 2.070 1.525 ;
        RECT  1.945 0.275 2.055 0.625 ;
        RECT  1.840 0.715 1.950 1.090 ;
        RECT  1.750 0.525 1.945 0.625 ;
        RECT  1.750 1.180 1.925 1.300 ;
        RECT  1.550 0.305 1.825 0.415 ;
        RECT  1.645 1.390 1.825 1.525 ;
        RECT  1.650 0.525 1.750 1.300 ;
        RECT  0.570 1.010 1.650 1.100 ;
        RECT  1.450 0.305 1.550 0.900 ;
        RECT  1.375 1.200 1.550 1.525 ;
        RECT  1.375 0.305 1.450 0.415 ;
        RECT  1.030 0.510 1.140 0.910 ;
        RECT  0.460 0.730 0.570 1.100 ;
        RECT  0.340 1.010 0.460 1.100 ;
        RECT  0.240 0.730 0.340 1.100 ;
        LAYER VIA1 ;
        RECT  2.480 1.415 2.580 1.515 ;
        RECT  2.450 0.750 2.550 0.850 ;
        RECT  2.210 1.190 2.310 1.290 ;
        RECT  1.910 1.415 2.010 1.515 ;
        RECT  1.450 0.750 1.550 0.850 ;
        RECT  1.450 1.290 1.550 1.390 ;
        LAYER M2 ;
        RECT  1.870 1.415 2.620 1.515 ;
        RECT  2.450 0.710 2.550 1.290 ;
        RECT  1.550 1.190 2.450 1.290 ;
        RECT  1.450 0.710 1.550 1.430 ;
    END
END GXOR2D2

MACRO HA1D0
    CLASS CORE ;
    FOREIGN HA1D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.480 3.150 1.290 ;
        RECT  3.025 0.480 3.050 0.695 ;
        RECT  3.025 1.045 3.050 1.290 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.275 0.175 0.485 ;
        RECT  0.150 1.280 0.175 1.490 ;
        RECT  0.050 0.275 0.150 1.490 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.1050 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.415 2.730 1.525 ;
        RECT  1.650 1.215 1.750 1.525 ;
        RECT  0.955 1.215 1.650 1.305 ;
        RECT  0.845 1.000 0.955 1.305 ;
        RECT  0.750 1.000 0.845 1.100 ;
        RECT  0.650 0.710 0.750 1.100 ;
        RECT  0.445 0.710 0.650 0.890 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0823 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 1.150 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.865 -0.165 3.200 0.165 ;
        RECT  2.755 -0.165 2.865 0.675 ;
        RECT  0.475 -0.165 2.755 0.165 ;
        RECT  0.305 -0.165 0.475 0.420 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.635 3.200 1.965 ;
        RECT  1.170 1.395 1.535 1.505 ;
        RECT  1.030 1.395 1.170 1.965 ;
        RECT  0.815 1.395 1.030 1.505 ;
        RECT  0.475 1.635 1.030 1.965 ;
        RECT  0.305 1.370 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.900 0.765 2.940 0.965 ;
        RECT  2.800 0.765 2.900 1.325 ;
        RECT  1.995 1.225 2.800 1.325 ;
        RECT  2.520 1.025 2.655 1.135 ;
        RECT  2.520 0.275 2.600 0.865 ;
        RECT  2.490 0.275 2.520 1.135 ;
        RECT  2.410 0.725 2.490 1.135 ;
        RECT  2.210 0.275 2.320 1.135 ;
        RECT  1.450 0.275 2.210 0.365 ;
        RECT  2.130 1.025 2.210 1.135 ;
        RECT  1.995 0.455 2.085 0.555 ;
        RECT  1.895 0.455 1.995 1.325 ;
        RECT  1.860 1.225 1.895 1.325 ;
        RECT  1.705 0.455 1.805 1.125 ;
        RECT  1.615 0.455 1.705 0.555 ;
        RECT  1.585 1.015 1.705 1.125 ;
        RECT  1.450 0.760 1.615 0.870 ;
        RECT  1.340 0.275 1.450 1.125 ;
        RECT  1.065 0.275 1.340 0.445 ;
        RECT  1.065 1.015 1.340 1.125 ;
        RECT  0.855 0.275 0.965 0.600 ;
        RECT  0.355 0.510 0.855 0.600 ;
        RECT  0.595 1.190 0.705 1.490 ;
        RECT  0.355 1.190 0.595 1.280 ;
        RECT  0.265 0.510 0.355 1.280 ;
        RECT  0.260 0.750 0.265 0.930 ;
    END
END HA1D0

MACRO HA1D1
    CLASS CORE ;
    FOREIGN HA1D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.225 0.275 3.350 1.500 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.275 0.175 0.675 ;
        RECT  0.150 1.045 0.175 1.505 ;
        RECT  0.050 0.275 0.150 1.505 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.1327 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.415 2.940 1.525 ;
        RECT  1.800 1.215 1.910 1.525 ;
        RECT  0.955 1.215 1.800 1.305 ;
        RECT  0.845 1.000 0.955 1.305 ;
        RECT  0.750 1.000 0.845 1.100 ;
        RECT  0.650 0.700 0.750 1.100 ;
        RECT  0.445 0.700 0.650 0.920 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1643 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.355 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.060 -0.165 3.400 0.165 ;
        RECT  2.950 -0.165 3.060 0.675 ;
        RECT  1.215 -0.165 2.950 0.165 ;
        RECT  1.105 -0.165 1.215 0.580 ;
        RECT  0.485 -0.165 1.105 0.165 ;
        RECT  0.295 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.635 3.400 1.965 ;
        RECT  1.420 1.395 1.610 1.965 ;
        RECT  1.005 1.635 1.420 1.965 ;
        RECT  0.815 1.395 1.005 1.965 ;
        RECT  0.485 1.635 0.815 1.965 ;
        RECT  0.295 1.395 0.485 1.965 ;
        RECT  0.000 1.635 0.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.100 0.775 3.135 0.955 ;
        RECT  3.000 0.775 3.100 1.325 ;
        RECT  2.195 1.225 3.000 1.325 ;
        RECT  2.720 1.025 2.840 1.135 ;
        RECT  2.720 0.275 2.790 0.865 ;
        RECT  2.680 0.275 2.720 1.135 ;
        RECT  2.610 0.725 2.680 1.135 ;
        RECT  2.410 0.275 2.520 1.135 ;
        RECT  1.555 0.275 2.410 0.365 ;
        RECT  2.320 1.025 2.410 1.135 ;
        RECT  2.195 0.455 2.275 0.555 ;
        RECT  2.095 0.455 2.195 1.325 ;
        RECT  2.020 1.225 2.095 1.325 ;
        RECT  1.905 0.455 2.005 1.125 ;
        RECT  1.825 0.455 1.905 0.555 ;
        RECT  1.755 1.015 1.905 1.125 ;
        RECT  1.555 0.720 1.815 0.910 ;
        RECT  1.445 0.275 1.555 1.125 ;
        RECT  1.325 0.275 1.445 0.445 ;
        RECT  1.065 1.015 1.445 1.125 ;
        RECT  0.815 0.275 0.985 0.610 ;
        RECT  0.355 0.500 0.815 0.610 ;
        RECT  0.595 1.215 0.705 1.495 ;
        RECT  0.355 1.215 0.595 1.305 ;
        RECT  0.265 0.500 0.355 1.305 ;
        RECT  0.260 0.750 0.265 0.930 ;
    END
END HA1D1

MACRO HA1D2
    CLASS CORE ;
    FOREIGN HA1D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.275 3.550 1.505 ;
        RECT  3.375 0.275 3.450 0.675 ;
        RECT  3.375 1.055 3.450 1.505 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.275 0.425 0.675 ;
        RECT  0.350 1.055 0.425 1.505 ;
        RECT  0.250 0.275 0.350 1.505 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.1334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.110 1.415 3.120 1.525 ;
        RECT  2.000 1.215 2.110 1.525 ;
        RECT  1.155 1.215 2.000 1.305 ;
        RECT  1.045 1.000 1.155 1.305 ;
        RECT  0.950 1.000 1.045 1.100 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.695 0.700 0.850 0.920 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1648 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.555 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.825 1.635 3.800 1.965 ;
        RECT  1.635 1.395 1.825 1.965 ;
        RECT  1.235 1.635 1.635 1.965 ;
        RECT  1.045 1.395 1.235 1.965 ;
        RECT  0.000 1.635 1.045 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.280 0.775 3.340 0.955 ;
        RECT  3.190 0.775 3.280 1.325 ;
        RECT  2.390 1.225 3.190 1.325 ;
        RECT  2.900 1.025 3.025 1.135 ;
        RECT  2.900 0.275 2.975 0.865 ;
        RECT  2.865 0.275 2.900 1.135 ;
        RECT  2.800 0.725 2.865 1.135 ;
        RECT  2.780 0.725 2.800 0.925 ;
        RECT  2.660 1.025 2.710 1.135 ;
        RECT  2.660 0.275 2.705 0.650 ;
        RECT  2.570 0.275 2.660 1.135 ;
        RECT  1.755 0.275 2.570 0.365 ;
        RECT  2.520 1.025 2.570 1.135 ;
        RECT  2.390 0.455 2.460 0.555 ;
        RECT  2.290 0.455 2.390 1.325 ;
        RECT  2.220 1.225 2.290 1.325 ;
        RECT  2.100 0.455 2.200 1.125 ;
        RECT  2.010 0.455 2.100 0.555 ;
        RECT  1.965 1.015 2.100 1.125 ;
        RECT  1.755 0.740 1.990 0.925 ;
        RECT  1.645 0.275 1.755 1.125 ;
        RECT  1.500 0.275 1.645 0.445 ;
        RECT  1.295 1.015 1.645 1.125 ;
        RECT  1.015 0.275 1.185 0.610 ;
        RECT  0.605 0.500 1.015 0.610 ;
        RECT  0.825 1.215 0.935 1.485 ;
        RECT  0.605 1.215 0.825 1.305 ;
        RECT  0.515 0.500 0.605 1.305 ;
        RECT  0.460 0.765 0.515 0.955 ;
    END
END HA1D2

MACRO HA1D4
    CLASS CORE ;
    FOREIGN HA1D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.300 5.550 0.670 ;
        RECT  5.450 1.100 5.550 1.470 ;
        RECT  5.150 0.300 5.450 1.470 ;
        RECT  4.825 0.300 5.150 0.670 ;
        RECT  4.825 1.100 5.150 1.470 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.300 0.940 0.670 ;
        RECT  0.650 1.100 0.940 1.470 ;
        RECT  0.350 0.300 0.650 1.470 ;
        RECT  0.250 0.300 0.350 0.670 ;
        RECT  0.250 1.100 0.350 1.470 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.1887 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.175 1.435 4.535 1.525 ;
        RECT  2.150 1.000 2.175 1.525 ;
        RECT  2.085 0.710 2.150 1.525 ;
        RECT  1.970 0.710 2.085 1.100 ;
        RECT  1.355 1.000 1.970 1.100 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.2755 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.710 2.705 0.890 ;
        RECT  2.250 0.510 2.350 0.890 ;
        RECT  1.755 0.510 2.250 0.610 ;
        RECT  1.650 0.510 1.755 0.890 ;
        RECT  1.535 0.785 1.650 0.890 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.825 0.300 5.050 0.670 ;
        RECT  4.825 1.100 5.050 1.470 ;
        RECT  0.750 0.300 0.940 0.670 ;
        RECT  0.750 1.100 0.940 1.470 ;
        RECT  4.715 0.800 4.960 0.900 ;
        RECT  4.615 0.800 4.715 1.345 ;
        RECT  3.905 1.255 4.615 1.345 ;
        RECT  4.365 0.275 4.475 1.165 ;
        RECT  4.335 0.745 4.365 1.165 ;
        RECT  4.285 0.745 4.335 0.915 ;
        RECT  4.160 0.275 4.220 0.650 ;
        RECT  4.160 0.995 4.220 1.165 ;
        RECT  4.065 0.275 4.160 1.165 ;
        RECT  2.925 0.275 4.065 0.365 ;
        RECT  3.905 0.455 3.975 0.570 ;
        RECT  3.805 0.455 3.905 1.345 ;
        RECT  3.615 0.455 3.715 1.250 ;
        RECT  3.035 0.455 3.615 0.555 ;
        RECT  3.045 1.140 3.615 1.250 ;
        RECT  2.925 0.790 3.470 0.900 ;
        RECT  2.825 0.275 2.925 1.280 ;
        RECT  2.295 0.275 2.825 0.420 ;
        RECT  2.285 1.160 2.825 1.280 ;
        RECT  1.140 1.215 1.975 1.335 ;
        RECT  0.870 0.790 1.050 0.910 ;
        RECT  1.140 0.310 1.735 0.420 ;
        RECT  1.050 0.310 1.140 1.335 ;
    END
END HA1D4

MACRO HCOSCIND1
    CLASS CORE ;
    FOREIGN HCOSCIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.275 5.950 1.490 ;
        RECT  5.815 0.275 5.850 0.675 ;
        RECT  5.815 1.045 5.850 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0659 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.710 4.550 0.905 ;
        END
    END CS
    PIN CO
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.275 0.175 0.675 ;
        RECT  0.150 1.045 0.175 1.490 ;
        RECT  0.050 0.275 0.150 1.490 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.700 3.950 0.900 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.2750 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.355 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.165 6.000 0.165 ;
        RECT  0.295 -0.165 0.485 0.405 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.635 6.000 1.965 ;
        RECT  5.490 1.510 5.660 1.965 ;
        RECT  3.915 1.635 5.490 1.965 ;
        RECT  3.745 1.370 3.915 1.965 ;
        RECT  2.185 1.635 3.745 1.965 ;
        RECT  2.015 1.415 2.185 1.965 ;
        RECT  0.970 1.635 2.015 1.965 ;
        RECT  0.970 1.395 1.595 1.505 ;
        RECT  0.830 1.395 0.970 1.965 ;
        RECT  0.305 1.395 0.830 1.505 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.765 5.760 0.955 ;
        RECT  5.605 0.765 5.705 1.400 ;
        RECT  4.895 1.310 5.605 1.400 ;
        RECT  5.315 0.455 5.425 1.175 ;
        RECT  5.180 0.825 5.315 0.935 ;
        RECT  5.070 1.025 5.205 1.115 ;
        RECT  5.070 0.275 5.165 0.735 ;
        RECT  5.055 0.275 5.070 1.115 ;
        RECT  3.375 0.275 5.055 0.365 ;
        RECT  4.980 0.645 5.055 1.115 ;
        RECT  4.870 0.455 4.935 0.565 ;
        RECT  4.870 1.165 4.895 1.400 ;
        RECT  4.765 0.455 4.870 1.400 ;
        RECT  4.160 0.455 4.675 0.565 ;
        RECT  4.160 1.205 4.675 1.315 ;
        RECT  4.050 0.455 4.160 1.490 ;
        RECT  4.020 0.455 4.050 0.565 ;
        RECT  3.555 0.475 3.745 0.585 ;
        RECT  3.555 1.090 3.745 1.230 ;
        RECT  3.465 0.475 3.555 1.525 ;
        RECT  3.310 1.435 3.465 1.525 ;
        RECT  3.285 0.275 3.375 1.295 ;
        RECT  3.120 1.385 3.310 1.525 ;
        RECT  2.605 1.205 3.285 1.295 ;
        RECT  3.085 0.410 3.195 1.115 ;
        RECT  2.365 1.435 3.120 1.525 ;
        RECT  2.945 0.695 3.085 0.865 ;
        RECT  2.855 1.025 2.975 1.115 ;
        RECT  2.855 0.475 2.945 0.585 ;
        RECT  2.765 0.275 2.855 1.115 ;
        RECT  1.555 0.275 2.765 0.365 ;
        RECT  2.605 0.475 2.675 0.585 ;
        RECT  2.505 0.475 2.605 1.295 ;
        RECT  1.950 0.475 2.415 0.585 ;
        RECT  1.950 1.015 2.385 1.125 ;
        RECT  2.275 1.215 2.365 1.525 ;
        RECT  0.955 1.215 2.275 1.305 ;
        RECT  1.850 0.475 1.950 1.125 ;
        RECT  1.760 0.475 1.850 0.585 ;
        RECT  1.700 1.015 1.850 1.125 ;
        RECT  1.555 0.720 1.760 0.910 ;
        RECT  1.445 0.275 1.555 1.125 ;
        RECT  1.260 0.275 1.445 0.445 ;
        RECT  1.075 1.015 1.445 1.125 ;
        RECT  0.940 0.500 0.975 0.610 ;
        RECT  0.845 1.000 0.955 1.305 ;
        RECT  0.820 0.275 0.940 0.610 ;
        RECT  0.580 1.000 0.845 1.100 ;
        RECT  0.355 0.500 0.820 0.610 ;
        RECT  0.355 1.195 0.745 1.305 ;
        RECT  0.450 0.700 0.580 1.100 ;
        RECT  0.265 0.500 0.355 1.305 ;
        RECT  0.240 0.765 0.265 0.955 ;
    END
END HCOSCIND1

MACRO HCOSCIND2
    CLASS CORE ;
    FOREIGN HCOSCIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.535 6.350 1.200 ;
        RECT  6.230 0.535 6.250 0.675 ;
        RECT  6.225 1.045 6.250 1.200 ;
        RECT  6.125 0.275 6.230 0.675 ;
        RECT  6.125 1.045 6.225 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0661 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.710 4.770 1.095 ;
        END
    END CS
    PIN CO
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.275 0.435 0.675 ;
        RECT  0.350 1.045 0.435 1.490 ;
        RECT  0.335 0.275 0.350 1.490 ;
        RECT  0.250 0.510 0.335 1.200 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.710 4.150 1.095 ;
        RECT  3.950 0.710 4.050 0.920 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.2750 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.555 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.490 -0.165 6.600 0.165 ;
        RECT  6.380 -0.165 6.490 0.445 ;
        RECT  5.970 -0.165 6.380 0.165 ;
        RECT  5.860 -0.165 5.970 0.675 ;
        RECT  0.745 -0.165 5.860 0.165 ;
        RECT  0.555 -0.165 0.745 0.405 ;
        RECT  0.185 -0.165 0.555 0.165 ;
        RECT  0.075 -0.165 0.185 0.445 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.490 1.635 6.600 1.965 ;
        RECT  6.380 1.315 6.490 1.965 ;
        RECT  5.945 1.635 6.380 1.965 ;
        RECT  5.775 1.490 5.945 1.965 ;
        RECT  4.175 1.635 5.775 1.965 ;
        RECT  4.005 1.425 4.175 1.965 ;
        RECT  2.445 1.635 4.005 1.965 ;
        RECT  2.275 1.415 2.445 1.965 ;
        RECT  1.170 1.635 2.275 1.965 ;
        RECT  1.170 1.395 1.845 1.500 ;
        RECT  1.030 1.395 1.170 1.965 ;
        RECT  0.555 1.395 1.030 1.500 ;
        RECT  0.185 1.635 1.030 1.965 ;
        RECT  0.075 1.355 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.000 0.810 6.140 0.910 ;
        RECT  5.900 0.810 6.000 1.400 ;
        RECT  5.155 1.310 5.900 1.400 ;
        RECT  5.575 0.455 5.685 1.175 ;
        RECT  5.440 0.825 5.575 0.935 ;
        RECT  5.330 1.025 5.465 1.115 ;
        RECT  5.330 0.275 5.425 0.735 ;
        RECT  5.315 0.275 5.330 1.115 ;
        RECT  3.635 0.275 5.315 0.365 ;
        RECT  5.240 0.645 5.315 1.115 ;
        RECT  5.130 0.455 5.195 0.565 ;
        RECT  5.130 1.165 5.155 1.400 ;
        RECT  5.025 0.455 5.130 1.400 ;
        RECT  4.420 0.455 4.935 0.565 ;
        RECT  4.420 1.205 4.935 1.315 ;
        RECT  4.310 0.455 4.420 1.490 ;
        RECT  4.280 0.455 4.310 0.565 ;
        RECT  3.815 0.475 3.985 0.585 ;
        RECT  3.815 1.065 3.950 1.255 ;
        RECT  3.725 0.475 3.815 1.525 ;
        RECT  3.570 1.435 3.725 1.525 ;
        RECT  3.545 0.275 3.635 1.295 ;
        RECT  3.380 1.385 3.570 1.525 ;
        RECT  2.865 1.205 3.545 1.295 ;
        RECT  3.345 0.410 3.455 1.115 ;
        RECT  2.625 1.435 3.380 1.525 ;
        RECT  3.205 0.695 3.345 0.865 ;
        RECT  3.115 1.025 3.235 1.115 ;
        RECT  3.115 0.475 3.205 0.585 ;
        RECT  3.025 0.275 3.115 1.115 ;
        RECT  1.815 0.275 3.025 0.365 ;
        RECT  2.865 0.475 2.935 0.585 ;
        RECT  2.765 0.475 2.865 1.295 ;
        RECT  2.210 0.475 2.675 0.585 ;
        RECT  2.210 1.015 2.645 1.125 ;
        RECT  2.535 1.215 2.625 1.525 ;
        RECT  1.225 1.215 2.535 1.305 ;
        RECT  2.110 0.475 2.210 1.125 ;
        RECT  2.020 0.475 2.110 0.585 ;
        RECT  1.960 1.015 2.110 1.125 ;
        RECT  1.815 0.720 2.020 0.910 ;
        RECT  1.705 0.275 1.815 1.125 ;
        RECT  1.520 0.275 1.705 0.445 ;
        RECT  1.335 1.015 1.705 1.125 ;
        RECT  1.080 0.275 1.235 0.610 ;
        RECT  1.115 1.000 1.225 1.305 ;
        RECT  0.840 1.000 1.115 1.100 ;
        RECT  0.615 0.500 1.080 0.610 ;
        RECT  0.615 1.215 1.005 1.305 ;
        RECT  0.710 0.700 0.840 1.100 ;
        RECT  0.525 0.500 0.615 1.305 ;
        RECT  0.500 0.765 0.525 0.955 ;
    END
END HCOSCIND2

MACRO HCOSCOND1
    CLASS CORE ;
    FOREIGN HCOSCOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.275 5.150 1.490 ;
        RECT  5.015 0.275 5.050 0.675 ;
        RECT  5.015 1.045 5.050 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0659 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.750 0.905 ;
        END
    END CS
    PIN CON
        ANTENNADIFFAREA 0.1620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.445 0.665 0.580 ;
        RECT  0.450 0.310 0.550 1.125 ;
        RECT  0.285 1.015 0.450 1.125 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.1012 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.665 1.385 2.855 1.525 ;
        RECT  2.035 1.435 2.665 1.525 ;
        RECT  1.945 1.215 2.035 1.525 ;
        RECT  0.170 1.215 1.945 1.305 ;
        RECT  0.050 0.710 0.170 1.305 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.2704 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.700 0.955 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.860 1.635 5.200 1.965 ;
        RECT  4.690 1.510 4.860 1.965 ;
        RECT  3.115 1.635 4.690 1.965 ;
        RECT  2.945 1.405 3.115 1.965 ;
        RECT  1.855 1.635 2.945 1.965 ;
        RECT  1.685 1.415 1.855 1.965 ;
        RECT  0.970 1.635 1.685 1.965 ;
        RECT  0.970 1.395 1.265 1.500 ;
        RECT  0.830 1.395 0.970 1.965 ;
        RECT  0.535 1.395 0.830 1.500 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.905 0.765 4.960 0.955 ;
        RECT  4.805 0.765 4.905 1.400 ;
        RECT  4.095 1.310 4.805 1.400 ;
        RECT  4.515 0.455 4.625 1.175 ;
        RECT  4.380 0.825 4.515 0.935 ;
        RECT  4.270 1.025 4.405 1.115 ;
        RECT  4.270 0.275 4.365 0.735 ;
        RECT  4.255 0.275 4.270 1.115 ;
        RECT  3.075 0.275 4.255 0.365 ;
        RECT  4.180 0.645 4.255 1.115 ;
        RECT  4.070 0.455 4.135 0.565 ;
        RECT  4.070 1.165 4.095 1.400 ;
        RECT  3.965 0.455 4.070 1.400 ;
        RECT  3.360 0.455 3.875 0.565 ;
        RECT  3.360 1.205 3.875 1.315 ;
        RECT  3.250 0.455 3.360 1.490 ;
        RECT  3.220 0.455 3.250 0.565 ;
        RECT  2.975 0.275 3.075 1.295 ;
        RECT  2.275 1.205 2.975 1.295 ;
        RECT  2.755 0.440 2.865 1.115 ;
        RECT  2.675 0.695 2.755 0.865 ;
        RECT  2.545 1.025 2.645 1.115 ;
        RECT  2.545 0.475 2.635 0.585 ;
        RECT  2.455 0.275 2.545 1.115 ;
        RECT  1.250 0.275 2.455 0.365 ;
        RECT  2.295 0.475 2.365 0.585 ;
        RECT  2.275 0.475 2.295 0.895 ;
        RECT  2.195 0.475 2.275 1.295 ;
        RECT  2.165 0.795 2.195 1.295 ;
        RECT  1.700 0.475 2.105 0.585 ;
        RECT  1.700 1.015 2.055 1.125 ;
        RECT  1.600 0.475 1.700 1.125 ;
        RECT  1.450 0.475 1.600 0.585 ;
        RECT  1.390 1.015 1.600 1.125 ;
        RECT  1.250 0.750 1.510 0.920 ;
        RECT  1.150 0.275 1.250 1.125 ;
        RECT  0.950 0.275 1.150 0.445 ;
        RECT  0.805 1.015 1.150 1.125 ;
    END
END HCOSCOND1

MACRO HCOSCOND2
    CLASS CORE ;
    FOREIGN HCOSCOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.665 0.545 5.750 1.200 ;
        RECT  5.650 0.275 5.665 1.490 ;
        RECT  5.555 0.275 5.650 0.690 ;
        RECT  5.555 1.045 5.650 1.490 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0659 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.710 4.350 0.905 ;
        END
    END CS
    PIN CON
        ANTENNADIFFAREA 0.2860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 1.015 1.025 1.125 ;
        RECT  0.555 0.310 0.775 0.435 ;
        RECT  0.445 0.310 0.555 1.125 ;
        RECT  0.315 1.015 0.445 1.125 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.1553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.205 1.385 3.395 1.525 ;
        RECT  2.575 1.435 3.205 1.525 ;
        RECT  2.485 1.215 2.575 1.525 ;
        RECT  1.250 1.215 2.485 1.305 ;
        RECT  1.150 0.735 1.250 1.305 ;
        RECT  1.050 0.735 1.150 0.905 ;
        RECT  0.170 1.215 1.150 1.305 ;
        RECT  0.050 0.710 0.170 1.305 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.3245 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.555 1.550 0.910 ;
        RECT  0.760 0.555 1.450 0.645 ;
        RECT  0.650 0.555 0.760 0.905 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.925 -0.165 6.000 0.165 ;
        RECT  5.815 -0.165 5.925 0.445 ;
        RECT  1.245 -0.165 5.815 0.165 ;
        RECT  1.125 -0.165 1.245 0.445 ;
        RECT  0.205 -0.165 1.125 0.165 ;
        RECT  0.095 -0.165 0.205 0.485 ;
        RECT  0.000 -0.165 0.095 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.925 1.635 6.000 1.965 ;
        RECT  5.815 1.355 5.925 1.965 ;
        RECT  5.400 1.635 5.815 1.965 ;
        RECT  5.230 1.510 5.400 1.965 ;
        RECT  3.655 1.635 5.230 1.965 ;
        RECT  3.485 1.425 3.655 1.965 ;
        RECT  2.395 1.635 3.485 1.965 ;
        RECT  2.225 1.415 2.395 1.965 ;
        RECT  1.370 1.635 2.225 1.965 ;
        RECT  1.370 1.395 1.815 1.500 ;
        RECT  1.230 1.395 1.370 1.965 ;
        RECT  0.560 1.395 1.230 1.500 ;
        RECT  0.000 1.635 1.230 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.445 0.810 5.560 0.910 ;
        RECT  5.345 0.810 5.445 1.400 ;
        RECT  4.635 1.310 5.345 1.400 ;
        RECT  5.055 0.455 5.165 1.175 ;
        RECT  4.920 0.825 5.055 0.935 ;
        RECT  4.810 1.025 4.945 1.115 ;
        RECT  4.810 0.275 4.905 0.735 ;
        RECT  4.795 0.275 4.810 1.115 ;
        RECT  3.615 0.275 4.795 0.365 ;
        RECT  4.720 0.645 4.795 1.115 ;
        RECT  4.610 0.455 4.675 0.565 ;
        RECT  4.610 1.165 4.635 1.400 ;
        RECT  4.505 0.455 4.610 1.400 ;
        RECT  3.900 0.455 4.415 0.565 ;
        RECT  3.900 1.205 4.415 1.315 ;
        RECT  3.790 0.455 3.900 1.490 ;
        RECT  3.760 0.455 3.790 0.565 ;
        RECT  3.515 0.275 3.615 1.295 ;
        RECT  2.815 1.205 3.515 1.295 ;
        RECT  3.295 0.440 3.405 1.115 ;
        RECT  3.215 0.695 3.295 0.865 ;
        RECT  3.085 1.025 3.185 1.115 ;
        RECT  3.085 0.475 3.175 0.585 ;
        RECT  2.995 0.275 3.085 1.115 ;
        RECT  1.790 0.275 2.995 0.365 ;
        RECT  2.835 0.475 2.905 0.585 ;
        RECT  2.815 0.475 2.835 0.895 ;
        RECT  2.735 0.475 2.815 1.295 ;
        RECT  2.705 0.795 2.735 1.295 ;
        RECT  2.370 0.475 2.645 0.585 ;
        RECT  2.370 1.015 2.595 1.125 ;
        RECT  2.270 0.475 2.370 1.125 ;
        RECT  1.880 0.475 2.270 0.585 ;
        RECT  1.930 1.015 2.270 1.125 ;
        RECT  1.790 0.765 2.110 0.905 ;
        RECT  1.690 0.275 1.790 1.125 ;
        RECT  1.355 0.275 1.690 0.420 ;
        RECT  1.355 1.015 1.690 1.125 ;
    END
END HCOSCOND2

MACRO HICIND1
    CLASS CORE ;
    FOREIGN HICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.275 3.750 1.490 ;
        RECT  3.615 0.275 3.650 0.675 ;
        RECT  3.615 1.045 3.650 1.490 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.275 0.175 0.675 ;
        RECT  0.150 1.045 0.175 1.490 ;
        RECT  0.050 0.275 0.150 1.490 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.1039 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.160 0.710 2.275 0.905 ;
        RECT  2.050 0.475 2.160 0.905 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.1648 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.355 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.165 3.800 0.165 ;
        RECT  0.295 -0.165 0.485 0.405 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.635 3.800 1.965 ;
        RECT  0.970 1.395 1.610 1.505 ;
        RECT  0.830 1.395 0.970 1.965 ;
        RECT  0.295 1.395 0.830 1.505 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.505 0.765 3.560 0.955 ;
        RECT  3.405 0.765 3.505 1.295 ;
        RECT  2.670 1.205 3.405 1.295 ;
        RECT  3.225 1.025 3.275 1.115 ;
        RECT  3.115 0.275 3.225 1.115 ;
        RECT  3.085 0.825 3.115 1.115 ;
        RECT  2.980 0.825 3.085 0.935 ;
        RECT  2.870 1.025 2.975 1.115 ;
        RECT  2.870 0.275 2.965 0.735 ;
        RECT  2.855 0.275 2.870 1.115 ;
        RECT  2.215 1.385 2.860 1.495 ;
        RECT  1.555 0.275 2.855 0.365 ;
        RECT  2.780 0.645 2.855 1.115 ;
        RECT  2.670 0.455 2.745 0.555 ;
        RECT  2.565 0.455 2.670 1.295 ;
        RECT  2.385 0.455 2.475 1.125 ;
        RECT  2.285 0.455 2.385 0.565 ;
        RECT  1.960 1.015 2.385 1.125 ;
        RECT  2.105 1.215 2.215 1.495 ;
        RECT  0.955 1.215 2.105 1.305 ;
        RECT  1.870 0.455 1.960 1.125 ;
        RECT  1.770 0.455 1.870 0.565 ;
        RECT  1.710 1.015 1.870 1.125 ;
        RECT  1.555 0.720 1.780 0.910 ;
        RECT  1.445 0.275 1.555 1.125 ;
        RECT  1.280 0.275 1.445 0.445 ;
        RECT  1.065 1.015 1.445 1.125 ;
        RECT  0.815 0.275 0.985 0.610 ;
        RECT  0.845 1.000 0.955 1.305 ;
        RECT  0.750 1.000 0.845 1.100 ;
        RECT  0.355 0.500 0.815 0.610 ;
        RECT  0.650 0.700 0.750 1.100 ;
        RECT  0.355 1.195 0.745 1.305 ;
        RECT  0.445 0.700 0.650 0.920 ;
        RECT  0.265 0.500 0.355 1.305 ;
        RECT  0.240 0.765 0.265 0.955 ;
    END
END HICIND1

MACRO HICIND2
    CLASS CORE ;
    FOREIGN HICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.275 3.950 1.490 ;
        RECT  3.775 0.275 3.850 0.675 ;
        RECT  3.775 1.055 3.850 1.490 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.295 0.485 0.410 ;
        RECT  0.150 1.390 0.485 1.490 ;
        RECT  0.050 0.295 0.150 1.490 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.1039 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.355 0.710 2.435 0.905 ;
        RECT  2.245 0.475 2.355 0.905 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.1648 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.555 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.570 1.635 4.200 1.965 ;
        RECT  1.570 1.395 1.800 1.505 ;
        RECT  1.430 1.395 1.570 1.965 ;
        RECT  1.045 1.395 1.430 1.505 ;
        RECT  0.000 1.635 1.430 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.685 0.765 3.740 0.955 ;
        RECT  3.585 0.765 3.685 1.295 ;
        RECT  2.805 1.205 3.585 1.295 ;
        RECT  3.375 1.025 3.425 1.115 ;
        RECT  3.265 0.485 3.375 1.115 ;
        RECT  3.235 0.725 3.265 1.115 ;
        RECT  3.180 0.725 3.235 0.905 ;
        RECT  3.080 0.275 3.175 0.445 ;
        RECT  3.080 0.995 3.120 1.115 ;
        RECT  2.980 0.275 3.080 1.115 ;
        RECT  2.795 1.385 2.995 1.525 ;
        RECT  1.755 0.275 2.980 0.365 ;
        RECT  2.915 0.995 2.980 1.115 ;
        RECT  2.805 0.455 2.890 0.565 ;
        RECT  2.705 0.455 2.805 1.295 ;
        RECT  2.085 1.415 2.795 1.525 ;
        RECT  2.525 0.455 2.615 1.125 ;
        RECT  2.445 0.455 2.525 0.565 ;
        RECT  2.155 1.015 2.525 1.125 ;
        RECT  2.045 0.455 2.155 1.125 ;
        RECT  1.975 1.215 2.085 1.525 ;
        RECT  1.940 0.455 2.045 0.555 ;
        RECT  1.880 1.015 2.045 1.125 ;
        RECT  1.155 1.215 1.975 1.305 ;
        RECT  1.755 0.720 1.950 0.910 ;
        RECT  1.645 0.275 1.755 1.125 ;
        RECT  1.450 0.275 1.645 0.445 ;
        RECT  1.305 1.015 1.645 1.125 ;
        RECT  0.985 0.275 1.155 0.610 ;
        RECT  1.045 0.990 1.155 1.305 ;
        RECT  0.950 0.990 1.045 1.090 ;
        RECT  0.500 0.500 0.985 0.610 ;
        RECT  0.850 0.700 0.950 1.090 ;
        RECT  0.825 1.200 0.935 1.470 ;
        RECT  0.650 0.700 0.850 0.920 ;
        RECT  0.500 1.200 0.825 1.290 ;
        RECT  0.390 0.500 0.500 1.290 ;
    END
END HICIND2

MACRO HICOND1
    CLASS CORE ;
    FOREIGN HICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.425 0.275 3.550 1.490 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.1660 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 0.275 0.750 0.690 ;
        RECT  0.150 0.555 0.605 0.690 ;
        RECT  0.150 1.180 0.525 1.290 ;
        RECT  0.050 0.555 0.150 1.290 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.1327 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 1.415 3.140 1.525 ;
        RECT  1.875 1.215 1.985 1.525 ;
        RECT  0.755 1.215 1.875 1.305 ;
        RECT  0.635 0.795 0.755 1.305 ;
        RECT  0.240 0.795 0.635 0.905 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.1648 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 1.155 0.900 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 -0.165 3.600 0.165 ;
        RECT  3.150 -0.165 3.260 0.660 ;
        RECT  0.215 -0.165 3.150 0.165 ;
        RECT  0.105 -0.165 0.215 0.445 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.635 3.600 1.965 ;
        RECT  1.170 1.395 1.360 1.965 ;
        RECT  0.765 1.635 1.170 1.965 ;
        RECT  0.595 1.395 0.765 1.965 ;
        RECT  0.000 1.635 0.595 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.300 0.765 3.335 0.955 ;
        RECT  3.200 0.765 3.300 1.325 ;
        RECT  2.395 1.225 3.200 1.325 ;
        RECT  2.920 1.025 3.040 1.135 ;
        RECT  2.920 0.275 2.990 0.865 ;
        RECT  2.880 0.275 2.920 1.135 ;
        RECT  2.810 0.725 2.880 1.135 ;
        RECT  2.610 0.275 2.720 1.135 ;
        RECT  1.355 0.275 2.610 0.365 ;
        RECT  2.520 1.025 2.610 1.135 ;
        RECT  2.395 0.455 2.485 0.555 ;
        RECT  2.295 0.455 2.395 1.325 ;
        RECT  2.215 1.225 2.295 1.325 ;
        RECT  2.105 0.455 2.205 1.115 ;
        RECT  1.540 0.455 2.105 0.565 ;
        RECT  1.480 1.015 2.105 1.115 ;
        RECT  1.355 0.720 1.550 0.910 ;
        RECT  1.245 0.275 1.355 1.125 ;
        RECT  1.050 0.275 1.245 0.445 ;
        RECT  0.845 1.015 1.245 1.125 ;
    END
END HICOND1

MACRO HICOND2
    CLASS CORE ;
    FOREIGN HICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.545 3.950 1.200 ;
        RECT  3.845 0.545 3.850 0.675 ;
        RECT  3.845 1.010 3.850 1.200 ;
        RECT  3.745 0.275 3.845 0.675 ;
        RECT  3.745 1.010 3.845 1.510 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.3020 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.215 1.035 1.305 ;
        RECT  0.150 0.310 0.765 0.420 ;
        RECT  0.050 0.310 0.150 1.305 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.1880 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.515 1.415 3.465 1.525 ;
        RECT  2.415 1.215 2.515 1.525 ;
        RECT  1.260 1.215 2.415 1.305 ;
        RECT  1.155 1.015 1.260 1.305 ;
        RECT  1.145 0.710 1.155 1.305 ;
        RECT  1.045 0.710 1.145 1.125 ;
        RECT  0.550 1.035 1.045 1.125 ;
        RECT  0.450 0.710 0.550 1.125 ;
        RECT  0.240 0.710 0.450 0.895 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.2191 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.510 1.555 0.925 ;
        RECT  0.750 0.510 1.445 0.610 ;
        RECT  0.650 0.510 0.750 0.925 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.110 -0.165 4.200 0.165 ;
        RECT  4.000 -0.165 4.110 0.465 ;
        RECT  3.585 -0.165 4.000 0.165 ;
        RECT  3.475 -0.165 3.585 0.680 ;
        RECT  1.285 -0.165 3.475 0.165 ;
        RECT  1.105 -0.165 1.285 0.405 ;
        RECT  0.000 -0.165 1.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.110 1.635 4.200 1.965 ;
        RECT  4.000 1.310 4.110 1.965 ;
        RECT  2.290 1.635 4.000 1.965 ;
        RECT  2.100 1.395 2.290 1.965 ;
        RECT  0.970 1.635 2.100 1.965 ;
        RECT  0.970 1.395 1.305 1.505 ;
        RECT  0.830 1.395 0.970 1.965 ;
        RECT  0.535 1.395 0.830 1.505 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.585 0.790 3.740 0.900 ;
        RECT  3.475 0.790 3.585 1.325 ;
        RECT  2.730 1.225 3.475 1.325 ;
        RECT  3.320 0.745 3.360 1.115 ;
        RECT  3.260 0.275 3.320 1.115 ;
        RECT  3.210 0.275 3.260 0.915 ;
        RECT  3.180 1.025 3.260 1.115 ;
        RECT  3.130 0.745 3.210 0.915 ;
        RECT  3.005 1.025 3.085 1.115 ;
        RECT  3.005 0.275 3.045 0.650 ;
        RECT  2.910 0.275 3.005 1.115 ;
        RECT  1.740 0.275 2.910 0.365 ;
        RECT  2.730 0.455 2.800 0.555 ;
        RECT  2.630 0.455 2.730 1.325 ;
        RECT  2.440 0.455 2.540 1.125 ;
        RECT  1.850 0.455 2.440 0.555 ;
        RECT  1.850 1.015 2.440 1.125 ;
        RECT  1.740 0.800 2.295 0.890 ;
        RECT  1.645 0.275 1.740 1.125 ;
        RECT  1.375 0.310 1.645 0.420 ;
        RECT  1.370 1.015 1.645 1.125 ;
    END
END HICOND2

MACRO IAO21D0
    CLASS CORE ;
    FOREIGN IAO21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0930 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.350 1.440 ;
        RECT  0.995 0.510 1.250 0.600 ;
        RECT  1.095 1.330 1.250 1.440 ;
        RECT  0.885 0.275 0.995 0.600 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.710 1.150 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 -0.165 1.400 0.165 ;
        RECT  1.215 0.300 1.305 0.400 ;
        RECT  1.105 -0.165 1.215 0.400 ;
        RECT  0.765 -0.165 1.105 0.165 ;
        RECT  0.595 -0.165 0.765 0.410 ;
        RECT  0.215 -0.165 0.595 0.165 ;
        RECT  0.105 -0.165 0.215 0.485 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.765 1.635 1.400 1.965 ;
        RECT  0.595 1.380 0.765 1.965 ;
        RECT  0.000 1.635 0.595 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 0.780 0.870 0.890 ;
        RECT  0.660 0.520 0.750 1.290 ;
        RECT  0.475 0.520 0.660 0.610 ;
        RECT  0.215 1.200 0.660 1.290 ;
        RECT  0.365 0.275 0.475 0.610 ;
        RECT  0.105 1.200 0.215 1.490 ;
    END
END IAO21D0

MACRO IAO21D1
    CLASS CORE ;
    FOREIGN IAO21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.350 1.310 ;
        RECT  0.995 0.510 1.250 0.600 ;
        RECT  1.095 1.200 1.250 1.310 ;
        RECT  0.885 0.370 0.995 0.600 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.710 1.150 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 -0.165 1.400 0.165 ;
        RECT  1.105 -0.165 1.285 0.400 ;
        RECT  0.765 -0.165 1.105 0.165 ;
        RECT  0.595 -0.165 0.765 0.410 ;
        RECT  0.215 -0.165 0.595 0.165 ;
        RECT  0.105 -0.165 0.215 0.485 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.765 1.635 1.400 1.965 ;
        RECT  0.595 1.380 0.765 1.965 ;
        RECT  0.000 1.635 0.595 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 0.780 0.870 0.890 ;
        RECT  0.660 0.520 0.750 1.290 ;
        RECT  0.475 0.520 0.660 0.610 ;
        RECT  0.215 1.200 0.660 1.290 ;
        RECT  0.365 0.275 0.475 0.610 ;
        RECT  0.105 1.200 0.215 1.490 ;
    END
END IAO21D1

MACRO IAO21D2
    CLASS CORE ;
    FOREIGN IAO21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.480 1.515 0.590 ;
        RECT  1.250 0.480 1.350 1.315 ;
        RECT  0.965 0.480 1.250 0.590 ;
        RECT  1.080 1.210 1.250 1.315 ;
        RECT  0.865 0.380 0.965 0.590 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.700 1.150 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.565 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.210 0.940 ;
        RECT  0.050 0.710 0.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.585 ;
        RECT  0.190 -0.165 1.615 0.165 ;
        RECT  0.080 -0.165 0.190 0.600 ;
        RECT  0.000 -0.165 0.080 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.635 1.800 1.965 ;
        RECT  0.575 1.395 0.750 1.965 ;
        RECT  0.000 1.635 0.575 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.560 0.730 1.670 1.495 ;
        RECT  0.970 1.405 1.560 1.495 ;
        RECT  0.895 1.210 0.970 1.495 ;
        RECT  0.880 0.780 0.895 1.495 ;
        RECT  0.805 0.780 0.880 1.305 ;
        RECT  0.775 0.780 0.805 0.890 ;
        RECT  0.205 1.210 0.805 1.305 ;
        RECT  0.685 0.480 0.775 0.890 ;
        RECT  0.305 0.480 0.685 0.590 ;
        RECT  0.095 1.210 0.205 1.420 ;
    END
END IAO21D2

MACRO IAO21D4
    CLASS CORE ;
    FOREIGN IAO21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.500 2.715 0.595 ;
        RECT  2.650 1.025 2.715 1.115 ;
        RECT  2.350 0.500 2.650 1.115 ;
        RECT  0.945 0.500 2.350 0.595 ;
        RECT  1.985 1.025 2.350 1.115 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0555 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.710 0.950 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.245 0.940 ;
        RECT  0.050 0.710 0.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.925 -0.165 3.000 0.165 ;
        RECT  2.815 -0.165 2.925 0.695 ;
        RECT  1.970 -0.165 2.815 0.165 ;
        RECT  1.970 0.305 2.455 0.410 ;
        RECT  1.830 -0.165 1.970 0.410 ;
        RECT  0.790 -0.165 1.830 0.165 ;
        RECT  1.205 0.305 1.830 0.410 ;
        RECT  0.650 -0.165 0.790 0.620 ;
        RECT  0.185 -0.165 0.650 0.165 ;
        RECT  0.075 -0.165 0.185 0.580 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.655 1.635 3.000 1.965 ;
        RECT  1.485 1.390 1.655 1.965 ;
        RECT  0.000 1.635 1.485 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.945 0.500 2.250 0.595 ;
        RECT  1.985 1.025 2.250 1.115 ;
        RECT  2.825 1.040 2.925 1.470 ;
        RECT  2.815 1.205 2.825 1.470 ;
        RECT  0.690 1.205 2.815 1.300 ;
        RECT  1.165 0.780 1.725 0.890 ;
        RECT  1.075 0.780 1.165 1.115 ;
        RECT  0.435 1.025 1.075 1.115 ;
        RECT  0.335 0.335 0.435 1.315 ;
        RECT  0.185 1.225 0.335 1.315 ;
        RECT  0.075 1.225 0.185 1.455 ;
    END
END IAO21D4

MACRO IAO22D0
    CLASS CORE ;
    FOREIGN IAO22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0830 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.330 1.255 0.440 ;
        RECT  1.050 0.330 1.150 1.090 ;
        RECT  0.950 1.000 1.050 1.090 ;
        RECT  0.840 1.000 0.950 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.530 0.710 1.650 0.940 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.365 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.260 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.490 ;
        RECT  0.945 -0.165 1.615 0.165 ;
        RECT  0.835 -0.165 0.945 0.470 ;
        RECT  0.190 -0.165 0.835 0.165 ;
        RECT  0.545 0.310 0.835 0.420 ;
        RECT  0.075 -0.165 0.190 0.485 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.495 1.635 1.800 1.965 ;
        RECT  1.325 1.385 1.495 1.965 ;
        RECT  0.190 1.635 1.325 1.965 ;
        RECT  0.070 1.280 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.615 1.200 1.725 1.490 ;
        RECT  1.205 1.200 1.615 1.295 ;
        RECT  1.095 1.200 1.205 1.490 ;
        RECT  0.750 0.780 0.960 0.890 ;
        RECT  0.660 0.530 0.750 1.440 ;
        RECT  0.445 0.530 0.660 0.620 ;
        RECT  0.525 1.330 0.660 1.440 ;
        RECT  0.335 0.275 0.445 0.620 ;
    END
END IAO22D0

MACRO IAO22D1
    CLASS CORE ;
    FOREIGN IAO22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.425 1.255 0.535 ;
        RECT  1.050 0.425 1.150 1.090 ;
        RECT  0.950 1.000 1.050 1.090 ;
        RECT  0.840 1.000 0.950 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.530 0.710 1.650 0.940 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.365 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.260 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.585 ;
        RECT  0.945 -0.165 1.615 0.165 ;
        RECT  0.840 -0.165 0.945 0.670 ;
        RECT  0.835 -0.165 0.840 0.420 ;
        RECT  0.190 -0.165 0.835 0.165 ;
        RECT  0.545 0.310 0.835 0.420 ;
        RECT  0.075 -0.165 0.190 0.485 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.495 1.635 1.800 1.965 ;
        RECT  1.325 1.385 1.495 1.965 ;
        RECT  0.190 1.635 1.325 1.965 ;
        RECT  0.070 1.280 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.615 1.200 1.725 1.410 ;
        RECT  1.045 1.200 1.615 1.295 ;
        RECT  0.750 0.780 0.960 0.890 ;
        RECT  0.660 0.530 0.750 1.440 ;
        RECT  0.445 0.530 0.660 0.620 ;
        RECT  0.525 1.330 0.660 1.440 ;
        RECT  0.335 0.275 0.445 0.620 ;
    END
END IAO22D1

MACRO IAO22D2
    CLASS CORE ;
    FOREIGN IAO22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.355 ;
        RECT  1.260 0.510 1.450 0.620 ;
        RECT  1.165 1.245 1.450 1.355 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0392 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.025 0.710 2.150 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0397 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.510 1.755 0.960 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.240 0.890 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.060 1.635 2.200 1.965 ;
        RECT  1.950 1.445 2.060 1.965 ;
        RECT  1.640 1.635 1.950 1.965 ;
        RECT  1.530 1.445 1.640 1.965 ;
        RECT  1.035 1.635 1.530 1.965 ;
        RECT  0.880 1.285 1.035 1.965 ;
        RECT  0.185 1.635 0.880 1.965 ;
        RECT  0.075 1.215 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.935 0.310 2.120 0.590 ;
        RECT  1.845 0.310 1.935 1.180 ;
        RECT  1.135 0.310 1.845 0.400 ;
        RECT  1.700 1.070 1.845 1.180 ;
        RECT  1.225 0.730 1.335 1.135 ;
        RECT  0.755 1.045 1.225 1.135 ;
        RECT  1.045 0.310 1.135 0.920 ;
        RECT  0.820 0.810 1.045 0.920 ;
        RECT  0.835 0.375 0.945 0.665 ;
        RECT  0.730 0.575 0.835 0.665 ;
        RECT  0.730 1.045 0.755 1.375 ;
        RECT  0.185 0.355 0.735 0.465 ;
        RECT  0.640 0.575 0.730 1.375 ;
        RECT  0.545 1.265 0.640 1.375 ;
        RECT  0.075 0.355 0.185 0.565 ;
    END
END IAO22D2

MACRO IAO22D4
    CLASS CORE ;
    FOREIGN IAO22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.015 2.815 1.120 ;
        RECT  2.675 0.275 2.785 0.695 ;
        RECT  2.650 0.520 2.675 0.695 ;
        RECT  2.350 0.520 2.650 1.120 ;
        RECT  2.105 0.520 2.350 0.630 ;
        RECT  2.125 1.015 2.350 1.120 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 0.710 3.550 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0395 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.030 0.710 3.150 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 1.150 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.560 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.045 -0.165 3.600 0.165 ;
        RECT  2.935 -0.165 3.045 0.585 ;
        RECT  2.370 -0.165 2.935 0.165 ;
        RECT  2.370 0.305 2.565 0.405 ;
        RECT  2.230 -0.165 2.370 0.405 ;
        RECT  0.770 -0.165 2.230 0.165 ;
        RECT  1.865 0.305 2.230 0.405 ;
        RECT  0.770 0.305 1.005 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.295 0.305 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 1.635 3.600 1.965 ;
        RECT  3.420 1.280 3.530 1.965 ;
        RECT  2.055 1.635 3.420 1.965 ;
        RECT  1.865 1.395 2.055 1.965 ;
        RECT  1.490 1.635 1.865 1.965 ;
        RECT  1.320 1.510 1.490 1.965 ;
        RECT  0.445 1.635 1.320 1.965 ;
        RECT  0.335 1.310 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 1.015 2.815 1.120 ;
        RECT  2.750 0.275 2.785 0.695 ;
        RECT  2.105 0.520 2.250 0.630 ;
        RECT  2.125 1.015 2.250 1.120 ;
        RECT  3.330 0.425 3.545 0.535 ;
        RECT  3.240 0.425 3.330 1.440 ;
        RECT  2.295 1.330 3.240 1.440 ;
        RECT  2.185 1.210 2.295 1.440 ;
        RECT  2.015 0.765 2.240 0.875 ;
        RECT  2.015 1.210 2.185 1.305 ;
        RECT  1.915 0.515 2.015 0.875 ;
        RECT  1.915 0.995 2.015 1.305 ;
        RECT  1.485 0.515 1.915 0.615 ;
        RECT  1.705 0.995 1.915 1.105 ;
        RECT  1.485 1.200 1.795 1.310 ;
        RECT  1.225 0.315 1.775 0.405 ;
        RECT  1.595 0.715 1.705 1.105 ;
        RECT  1.385 0.515 1.485 1.420 ;
        RECT  1.325 0.515 1.385 0.615 ;
        RECT  0.805 1.310 1.385 1.420 ;
        RECT  0.705 1.040 1.275 1.150 ;
        RECT  1.115 0.315 1.225 0.600 ;
        RECT  0.185 0.500 1.115 0.600 ;
        RECT  0.595 1.040 0.705 1.470 ;
        RECT  0.185 1.040 0.595 1.150 ;
        RECT  0.075 0.355 0.185 0.600 ;
        RECT  0.075 1.040 0.185 1.470 ;
    END
END IAO22D4

MACRO IIND4D0
    CLASS CORE ;
    FOREIGN IIND4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1380 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.275 1.405 0.485 ;
        RECT  1.250 0.275 1.350 1.160 ;
        RECT  1.225 1.050 1.250 1.160 ;
        RECT  1.115 1.050 1.225 1.490 ;
        RECT  0.705 1.050 1.115 1.160 ;
        RECT  0.595 1.050 0.705 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.780 0.830 0.890 ;
        RECT  0.650 0.510 0.750 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.890 ;
        RECT  0.920 0.780 1.050 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 1.950 1.090 ;
        RECT  1.810 0.710 1.850 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.695 -0.165 2.000 0.165 ;
        RECT  1.515 -0.165 1.695 0.420 ;
        RECT  0.475 -0.165 1.515 0.165 ;
        RECT  0.305 -0.165 0.475 0.420 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 1.635 2.000 1.965 ;
        RECT  1.375 1.270 1.485 1.965 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.835 1.270 0.965 1.965 ;
        RECT  0.475 1.635 0.835 1.965 ;
        RECT  0.305 1.380 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.815 0.285 1.925 0.600 ;
        RECT  1.695 0.510 1.815 0.600 ;
        RECT  1.695 1.330 1.795 1.440 ;
        RECT  1.585 0.510 1.695 1.440 ;
        RECT  1.440 0.785 1.585 0.890 ;
        RECT  0.390 0.780 0.560 0.890 ;
        RECT  0.300 0.510 0.390 1.290 ;
        RECT  0.185 0.510 0.300 0.600 ;
        RECT  0.185 1.200 0.300 1.290 ;
        RECT  0.075 0.275 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.490 ;
    END
END IIND4D0

MACRO IIND4D1
    CLASS CORE ;
    FOREIGN IIND4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.405 1.405 0.615 ;
        RECT  1.250 0.405 1.350 1.160 ;
        RECT  1.225 1.050 1.250 1.160 ;
        RECT  1.115 1.050 1.225 1.490 ;
        RECT  0.705 1.050 1.115 1.160 ;
        RECT  0.595 1.050 0.705 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.780 0.830 0.890 ;
        RECT  0.650 0.510 0.750 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.890 ;
        RECT  0.920 0.780 1.050 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 1.950 1.090 ;
        RECT  1.810 0.710 1.850 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.635 -0.165 2.000 0.165 ;
        RECT  1.635 0.310 1.705 0.420 ;
        RECT  1.515 -0.165 1.635 0.420 ;
        RECT  0.405 -0.165 1.515 0.165 ;
        RECT  0.405 0.310 0.495 0.420 ;
        RECT  0.295 -0.165 0.405 0.420 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 1.635 2.000 1.965 ;
        RECT  1.375 1.270 1.485 1.965 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.835 1.270 0.965 1.965 ;
        RECT  0.405 1.635 0.835 1.965 ;
        RECT  0.405 1.380 0.495 1.490 ;
        RECT  0.295 1.380 0.405 1.965 ;
        RECT  0.000 1.635 0.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.815 0.285 1.925 0.600 ;
        RECT  1.695 0.510 1.815 0.600 ;
        RECT  1.695 1.330 1.795 1.440 ;
        RECT  1.585 0.510 1.695 1.440 ;
        RECT  1.440 0.785 1.585 0.890 ;
        RECT  0.390 0.780 0.560 0.890 ;
        RECT  0.300 0.510 0.390 1.290 ;
        RECT  0.185 0.510 0.300 0.600 ;
        RECT  0.185 1.200 0.300 1.290 ;
        RECT  0.075 0.275 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.490 ;
    END
END IIND4D1

MACRO IIND4D2
    CLASS CORE ;
    FOREIGN IIND4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4940 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 1.010 3.065 1.130 ;
        RECT  1.155 0.510 1.270 0.630 ;
        RECT  1.050 0.510 1.155 1.130 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.560 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.790 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.065 -0.165 3.400 0.165 ;
        RECT  2.895 -0.165 3.065 0.405 ;
        RECT  0.475 -0.165 2.895 0.165 ;
        RECT  0.305 -0.165 0.475 0.420 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.325 1.635 3.400 1.965 ;
        RECT  3.155 1.400 3.325 1.965 ;
        RECT  2.805 1.635 3.155 1.965 ;
        RECT  2.635 1.400 2.805 1.965 ;
        RECT  2.185 1.635 2.635 1.965 ;
        RECT  2.185 1.400 2.310 1.515 ;
        RECT  2.015 1.400 2.185 1.965 ;
        RECT  1.835 1.400 2.015 1.515 ;
        RECT  1.505 1.635 2.015 1.965 ;
        RECT  1.335 1.400 1.505 1.965 ;
        RECT  0.985 1.635 1.335 1.965 ;
        RECT  0.815 1.400 0.985 1.965 ;
        RECT  0.475 1.635 0.815 1.965 ;
        RECT  0.305 1.400 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.345 3.295 0.600 ;
        RECT  3.175 0.775 3.285 1.310 ;
        RECT  2.775 0.500 3.185 0.600 ;
        RECT  2.880 0.775 3.175 0.890 ;
        RECT  0.350 1.220 3.175 1.310 ;
        RECT  2.665 0.310 2.775 0.600 ;
        RECT  2.115 0.310 2.665 0.410 ;
        RECT  1.575 0.520 2.555 0.620 ;
        RECT  0.950 0.310 2.025 0.410 ;
        RECT  0.750 0.770 0.960 0.900 ;
        RECT  0.840 0.310 0.950 0.590 ;
        RECT  0.640 0.295 0.750 1.130 ;
        RECT  0.565 0.295 0.640 0.405 ;
        RECT  0.545 1.020 0.640 1.130 ;
        RECT  0.260 0.510 0.350 1.310 ;
        RECT  0.185 0.510 0.260 0.600 ;
        RECT  0.185 1.220 0.260 1.310 ;
        RECT  0.075 0.375 0.185 0.600 ;
        RECT  0.075 1.220 0.185 1.420 ;
    END
END IIND4D2

MACRO IIND4D4
    CLASS CORE ;
    FOREIGN IIND4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.655 1.130 5.715 1.300 ;
        RECT  5.350 0.500 5.655 1.300 ;
        RECT  4.985 0.500 5.350 0.620 ;
        RECT  1.520 1.200 5.350 1.300 ;
        RECT  1.420 1.200 1.520 1.460 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.780 3.350 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.780 4.350 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.680 0.190 0.940 ;
        RECT  0.050 0.680 0.150 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.165 6.000 0.165 ;
        RECT  1.770 0.300 2.295 0.410 ;
        RECT  1.630 -0.165 1.770 0.410 ;
        RECT  0.705 -0.165 1.630 0.165 ;
        RECT  1.075 0.300 1.630 0.410 ;
        RECT  0.595 -0.165 0.705 0.560 ;
        RECT  0.185 -0.165 0.595 0.165 ;
        RECT  0.075 -0.165 0.185 0.560 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.925 1.635 6.000 1.965 ;
        RECT  5.815 1.040 5.925 1.965 ;
        RECT  5.170 1.635 5.815 1.965 ;
        RECT  5.170 1.390 5.455 1.500 ;
        RECT  5.030 1.390 5.170 1.965 ;
        RECT  4.465 1.390 5.030 1.500 ;
        RECT  3.570 1.635 5.030 1.965 ;
        RECT  3.570 1.390 4.155 1.500 ;
        RECT  3.430 1.390 3.570 1.965 ;
        RECT  2.905 1.390 3.430 1.500 ;
        RECT  2.170 1.635 3.430 1.965 ;
        RECT  2.170 1.390 2.595 1.500 ;
        RECT  2.030 1.390 2.170 1.965 ;
        RECT  1.630 1.390 2.030 1.500 ;
        RECT  0.970 1.635 2.030 1.965 ;
        RECT  0.970 1.390 1.310 1.495 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.555 1.390 0.830 1.495 ;
        RECT  0.185 1.635 0.830 1.965 ;
        RECT  0.075 1.240 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.985 0.500 5.250 0.620 ;
        RECT  1.520 1.200 5.250 1.300 ;
        RECT  1.420 1.200 1.520 1.460 ;
        RECT  5.815 0.305 5.925 0.585 ;
        RECT  3.695 0.305 5.815 0.410 ;
        RECT  5.045 0.730 5.155 1.090 ;
        RECT  1.330 1.000 5.045 1.090 ;
        RECT  3.585 0.500 4.675 0.600 ;
        RECT  3.475 0.305 3.585 0.600 ;
        RECT  2.405 0.305 3.475 0.410 ;
        RECT  1.325 0.500 3.365 0.600 ;
        RECT  1.130 0.780 2.070 0.890 ;
        RECT  1.240 1.000 1.330 1.300 ;
        RECT  0.445 1.210 1.240 1.300 ;
        RECT  1.040 0.510 1.130 1.120 ;
        RECT  0.965 0.510 1.040 0.600 ;
        RECT  0.805 1.015 1.040 1.120 ;
        RECT  0.855 0.350 0.965 0.600 ;
        RECT  0.335 0.350 0.445 1.475 ;
    END
END IIND4D4

MACRO IINR4D0
    CLASS CORE ;
    FOREIGN IINR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1510 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 0.275 1.310 0.470 ;
        RECT  0.750 0.380 1.200 0.470 ;
        RECT  0.625 0.275 0.750 1.130 ;
        RECT  0.500 1.020 0.625 1.130 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.710 1.550 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.710 1.215 0.920 ;
        RECT  1.050 0.710 1.150 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.710 1.950 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 -0.165 2.000 0.165 ;
        RECT  1.535 -0.165 1.645 0.420 ;
        RECT  1.060 -0.165 1.535 0.165 ;
        RECT  1.435 0.310 1.535 0.420 ;
        RECT  0.860 -0.165 1.060 0.290 ;
        RECT  0.405 -0.165 0.860 0.165 ;
        RECT  0.405 0.310 0.505 0.420 ;
        RECT  0.295 -0.165 0.405 0.420 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.635 2.000 1.965 ;
        RECT  1.170 1.390 1.640 1.500 ;
        RECT  1.030 1.390 1.170 1.965 ;
        RECT  0.295 1.390 1.030 1.500 ;
        RECT  0.000 1.635 1.030 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.740 1.200 1.930 1.300 ;
        RECT  1.770 0.275 1.880 0.600 ;
        RECT  1.740 0.510 1.770 0.600 ;
        RECT  1.640 0.510 1.740 1.300 ;
        RECT  0.960 1.200 1.640 1.300 ;
        RECT  0.860 0.560 0.960 1.300 ;
        RECT  0.370 0.735 0.535 0.905 ;
        RECT  0.280 0.510 0.370 1.290 ;
        RECT  0.185 0.510 0.280 0.600 ;
        RECT  0.185 1.200 0.280 1.290 ;
        RECT  0.075 0.275 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.480 ;
    END
END IINR4D0

MACRO IINR4D1
    CLASS CORE ;
    FOREIGN IINR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 0.285 1.900 0.610 ;
        RECT  1.150 0.500 1.790 0.610 ;
        RECT  1.150 1.185 1.550 1.295 ;
        RECT  1.050 0.500 1.150 1.295 ;
        RECT  0.055 0.500 1.050 0.610 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0753 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.750 1.090 ;
        RECT  0.620 0.710 0.650 0.940 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0754 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.170 0.710 0.250 0.940 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 2.350 0.890 ;
        RECT  2.200 0.700 2.250 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.700 2.570 0.910 ;
        RECT  2.450 0.510 2.550 0.910 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.165 2.800 0.165 ;
        RECT  2.430 0.295 2.490 0.400 ;
        RECT  2.320 -0.165 2.430 0.400 ;
        RECT  1.170 -0.165 2.320 0.165 ;
        RECT  1.170 0.305 1.680 0.410 ;
        RECT  1.030 -0.165 1.170 0.410 ;
        RECT  0.000 -0.165 1.030 0.165 ;
        RECT  0.330 0.305 1.030 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.635 2.800 1.965 ;
        RECT  2.370 1.405 2.560 1.965 ;
        RECT  0.685 1.635 2.370 1.965 ;
        RECT  0.575 1.390 0.685 1.965 ;
        RECT  0.485 1.390 0.575 1.495 ;
        RECT  0.000 1.635 0.575 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.660 0.295 2.750 1.295 ;
        RECT  2.580 0.295 2.660 0.400 ;
        RECT  2.615 1.025 2.660 1.295 ;
        RECT  1.750 1.205 2.615 1.295 ;
        RECT  2.090 1.010 2.275 1.115 ;
        RECT  2.090 0.295 2.230 0.400 ;
        RECT  2.000 0.295 2.090 1.115 ;
        RECT  0.885 1.385 2.015 1.485 ;
        RECT  1.860 0.750 2.000 0.920 ;
        RECT  1.660 0.775 1.750 1.295 ;
        RECT  1.360 0.775 1.660 0.890 ;
        RECT  0.795 1.210 0.885 1.485 ;
        RECT  0.185 1.210 0.795 1.300 ;
        RECT  0.075 1.210 0.185 1.415 ;
    END
END IINR4D1

MACRO IINR4D2
    CLASS CORE ;
    FOREIGN IINR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.155 1.155 4.840 1.265 ;
        RECT  4.155 0.480 4.570 0.590 ;
        RECT  4.045 0.480 4.155 1.265 ;
        RECT  3.030 0.480 4.045 0.590 ;
        RECT  2.920 0.390 3.030 0.590 ;
        RECT  1.180 0.390 2.920 0.485 ;
        RECT  1.080 0.300 1.180 0.485 ;
        RECT  0.895 0.300 1.080 0.410 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1719 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.770 1.555 1.105 ;
        RECT  0.650 0.770 1.445 0.900 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1722 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.770 2.555 0.900 ;
        RECT  2.050 0.770 2.350 1.105 ;
        RECT  1.845 0.770 2.050 0.900 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.255 0.930 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.420 0.710 5.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.170 -0.165 5.600 0.165 ;
        RECT  5.170 0.310 5.315 0.420 ;
        RECT  5.030 -0.165 5.170 0.420 ;
        RECT  4.790 -0.165 5.030 0.165 ;
        RECT  4.680 -0.165 4.790 0.685 ;
        RECT  3.970 -0.165 4.680 0.165 ;
        RECT  3.970 0.275 4.270 0.370 ;
        RECT  3.830 -0.165 3.970 0.370 ;
        RECT  3.010 -0.165 3.830 0.165 ;
        RECT  3.430 0.275 3.830 0.370 ;
        RECT  2.800 -0.165 3.010 0.300 ;
        RECT  2.600 -0.165 2.800 0.165 ;
        RECT  2.390 -0.165 2.600 0.300 ;
        RECT  1.920 -0.165 2.390 0.165 ;
        RECT  1.710 -0.165 1.920 0.300 ;
        RECT  1.500 -0.165 1.710 0.165 ;
        RECT  1.290 -0.165 1.500 0.300 ;
        RECT  0.570 -0.165 1.290 0.165 ;
        RECT  0.570 0.300 0.785 0.410 ;
        RECT  0.430 -0.165 0.570 0.410 ;
        RECT  0.000 -0.165 0.430 0.165 ;
        RECT  0.295 0.300 0.430 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.965 1.635 5.600 1.965 ;
        RECT  0.855 1.290 0.965 1.965 ;
        RECT  0.405 1.635 0.855 1.965 ;
        RECT  0.405 1.395 0.485 1.495 ;
        RECT  0.295 1.395 0.405 1.965 ;
        RECT  0.000 1.635 0.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.415 0.330 5.525 0.600 ;
        RECT  5.415 1.240 5.525 1.500 ;
        RECT  5.310 0.510 5.415 0.600 ;
        RECT  5.310 1.240 5.415 1.350 ;
        RECT  5.200 0.510 5.310 1.350 ;
        RECT  4.275 0.775 5.200 0.885 ;
        RECT  4.940 1.035 5.050 1.485 ;
        RECT  2.865 1.375 4.940 1.485 ;
        RECT  2.755 1.035 3.835 1.145 ;
        RECT  2.800 0.800 3.555 0.890 ;
        RECT  2.690 0.575 2.800 0.890 ;
        RECT  2.645 1.035 2.755 1.505 ;
        RECT  0.970 0.575 2.690 0.670 ;
        RECT  1.555 1.395 2.645 1.505 ;
        RECT  1.225 1.195 2.535 1.285 ;
        RECT  1.115 1.050 1.225 1.500 ;
        RECT  0.705 1.050 1.115 1.160 ;
        RECT  0.870 0.500 0.970 0.670 ;
        RECT  0.445 0.500 0.870 0.590 ;
        RECT  0.595 1.050 0.705 1.500 ;
        RECT  0.355 0.500 0.445 1.305 ;
        RECT  0.185 0.500 0.355 0.590 ;
        RECT  0.185 1.215 0.355 1.305 ;
        RECT  0.075 0.380 0.185 0.590 ;
        RECT  0.075 1.215 0.185 1.460 ;
    END
END IINR4D2

MACRO IINR4D4
    CLASS CORE ;
    FOREIGN IINR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 1.010 7.335 1.180 ;
        RECT  6.930 0.275 7.060 0.475 ;
        RECT  6.490 0.385 6.930 0.475 ;
        RECT  6.450 0.275 6.490 0.475 ;
        RECT  6.360 0.275 6.450 1.180 ;
        RECT  6.105 0.385 6.360 1.180 ;
        RECT  5.470 0.385 6.105 0.475 ;
        RECT  5.340 0.275 5.470 0.475 ;
        RECT  4.900 0.385 5.340 0.475 ;
        RECT  4.770 0.275 4.900 0.475 ;
        RECT  3.680 0.385 4.770 0.475 ;
        RECT  3.550 0.275 3.680 0.475 ;
        RECT  3.110 0.385 3.550 0.475 ;
        RECT  2.980 0.275 3.110 0.475 ;
        RECT  2.070 0.385 2.980 0.475 ;
        RECT  1.940 0.275 2.070 0.475 ;
        RECT  1.500 0.385 1.940 0.475 ;
        RECT  1.370 0.275 1.500 0.475 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2984 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.565 1.710 0.675 ;
        RECT  0.850 0.565 0.955 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2971 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 0.565 3.710 0.675 ;
        RECT  2.045 0.565 2.155 0.900 ;
        RECT  1.845 0.710 2.045 0.900 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.180 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.200 0.680 8.350 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.325 -0.165 8.400 0.165 ;
        RECT  8.215 -0.165 8.325 0.560 ;
        RECT  7.805 -0.165 8.215 0.165 ;
        RECT  7.695 -0.165 7.805 0.475 ;
        RECT  7.375 -0.165 7.695 0.165 ;
        RECT  7.245 -0.165 7.375 0.445 ;
        RECT  6.815 -0.165 7.245 0.165 ;
        RECT  6.605 -0.165 6.815 0.295 ;
        RECT  6.215 -0.165 6.605 0.165 ;
        RECT  6.005 -0.165 6.215 0.295 ;
        RECT  5.825 -0.165 6.005 0.165 ;
        RECT  5.615 -0.165 5.825 0.295 ;
        RECT  5.225 -0.165 5.615 0.165 ;
        RECT  5.020 -0.165 5.225 0.295 ;
        RECT  4.625 -0.165 5.020 0.165 ;
        RECT  4.415 -0.165 4.625 0.295 ;
        RECT  4.035 -0.165 4.415 0.165 ;
        RECT  3.825 -0.165 4.035 0.295 ;
        RECT  3.435 -0.165 3.825 0.165 ;
        RECT  3.225 -0.165 3.435 0.295 ;
        RECT  2.835 -0.165 3.225 0.165 ;
        RECT  2.625 -0.165 2.835 0.295 ;
        RECT  2.425 -0.165 2.625 0.165 ;
        RECT  2.215 -0.165 2.425 0.295 ;
        RECT  1.825 -0.165 2.215 0.165 ;
        RECT  1.615 -0.165 1.825 0.295 ;
        RECT  1.185 -0.165 1.615 0.165 ;
        RECT  1.055 -0.165 1.185 0.350 ;
        RECT  0.740 -0.165 1.055 0.165 ;
        RECT  0.610 -0.165 0.740 0.355 ;
        RECT  0.185 -0.165 0.610 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.325 1.635 8.400 1.965 ;
        RECT  8.215 1.260 8.325 1.965 ;
        RECT  7.815 1.635 8.215 1.965 ;
        RECT  7.685 0.980 7.815 1.965 ;
        RECT  1.805 1.635 7.685 1.965 ;
        RECT  1.635 1.460 1.805 1.965 ;
        RECT  1.235 1.635 1.635 1.965 ;
        RECT  1.065 1.460 1.235 1.965 ;
        RECT  0.185 1.635 1.065 1.965 ;
        RECT  0.075 1.260 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.550 1.010 7.335 1.180 ;
        RECT  6.930 0.275 7.060 0.475 ;
        RECT  6.550 0.385 6.930 0.475 ;
        RECT  5.470 0.385 6.050 0.475 ;
        RECT  5.340 0.275 5.470 0.475 ;
        RECT  4.900 0.385 5.340 0.475 ;
        RECT  4.770 0.275 4.900 0.475 ;
        RECT  3.680 0.385 4.770 0.475 ;
        RECT  3.550 0.275 3.680 0.475 ;
        RECT  3.110 0.385 3.550 0.475 ;
        RECT  2.980 0.275 3.110 0.475 ;
        RECT  2.070 0.385 2.980 0.475 ;
        RECT  1.940 0.275 2.070 0.475 ;
        RECT  1.500 0.385 1.940 0.475 ;
        RECT  1.370 0.275 1.500 0.475 ;
        RECT  7.960 0.350 8.065 1.470 ;
        RECT  7.955 0.350 7.960 0.675 ;
        RECT  6.600 0.565 7.955 0.675 ;
        RECT  7.435 0.980 7.545 1.445 ;
        RECT  5.985 1.335 7.435 1.445 ;
        RECT  5.875 0.865 5.985 1.445 ;
        RECT  5.465 1.335 5.875 1.445 ;
        RECT  5.615 0.775 5.725 1.225 ;
        RECT  5.205 0.775 5.615 0.895 ;
        RECT  5.355 0.995 5.465 1.445 ;
        RECT  4.335 0.565 5.410 0.665 ;
        RECT  4.945 1.335 5.355 1.445 ;
        RECT  5.095 0.775 5.205 1.225 ;
        RECT  4.735 0.775 5.095 0.885 ;
        RECT  4.835 0.995 4.945 1.445 ;
        RECT  4.275 1.335 4.835 1.445 ;
        RECT  4.625 0.775 4.735 1.140 ;
        RECT  2.705 1.030 4.625 1.140 ;
        RECT  4.205 0.565 4.335 0.915 ;
        RECT  2.585 0.785 4.205 0.915 ;
        RECT  4.055 1.240 4.165 1.510 ;
        RECT  0.770 1.240 4.055 1.350 ;
        RECT  2.465 0.785 2.585 1.140 ;
        RECT  0.445 1.010 2.465 1.140 ;
        RECT  0.335 0.375 0.445 1.500 ;
    END
END IINR4D4

MACRO IND2D0
    CLASS CORE ;
    FOREIGN IND2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.310 1.150 1.290 ;
        RECT  0.890 0.310 1.050 0.420 ;
        RECT  0.795 1.200 1.050 1.290 ;
        RECT  0.685 1.200 0.795 1.500 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0267 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.960 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0267 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.165 1.200 0.165 ;
        RECT  0.485 0.310 0.585 0.420 ;
        RECT  0.375 -0.165 0.485 0.420 ;
        RECT  0.000 -0.165 0.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.105 1.635 1.200 1.965 ;
        RECT  0.995 1.400 1.105 1.965 ;
        RECT  0.895 1.400 0.995 1.510 ;
        RECT  0.485 1.635 0.995 1.965 ;
        RECT  0.485 1.380 0.585 1.490 ;
        RECT  0.375 1.380 0.485 1.965 ;
        RECT  0.000 1.635 0.375 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.575 0.750 0.680 0.920 ;
        RECT  0.470 0.530 0.575 1.270 ;
        RECT  0.275 0.530 0.470 0.620 ;
        RECT  0.275 1.180 0.470 1.270 ;
        RECT  0.165 0.275 0.275 0.620 ;
        RECT  0.165 1.180 0.275 1.480 ;
    END
END IND2D0

MACRO IND2D1
    CLASS CORE ;
    FOREIGN IND2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.425 1.150 1.290 ;
        RECT  0.850 0.425 1.050 0.535 ;
        RECT  0.795 1.200 1.050 1.290 ;
        RECT  0.685 1.200 0.795 1.410 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.960 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 -0.165 1.200 0.165 ;
        RECT  0.495 0.310 0.585 0.420 ;
        RECT  0.385 -0.165 0.495 0.420 ;
        RECT  0.000 -0.165 0.385 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 1.635 1.200 1.965 ;
        RECT  1.015 1.400 1.105 1.500 ;
        RECT  0.905 1.400 1.015 1.965 ;
        RECT  0.485 1.635 0.905 1.965 ;
        RECT  0.485 1.380 0.585 1.490 ;
        RECT  0.375 1.380 0.485 1.965 ;
        RECT  0.000 1.635 0.375 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.575 0.750 0.680 0.920 ;
        RECT  0.485 0.530 0.575 1.270 ;
        RECT  0.275 0.530 0.485 0.620 ;
        RECT  0.275 1.180 0.485 1.270 ;
        RECT  0.165 0.275 0.275 0.620 ;
        RECT  0.165 1.180 0.275 1.480 ;
    END
END IND2D1

MACRO IND2D2
    CLASS CORE ;
    FOREIGN IND2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.050 1.255 1.480 ;
        RECT  1.145 0.510 1.150 1.480 ;
        RECT  1.050 0.510 1.145 1.285 ;
        RECT  0.840 0.510 1.050 0.620 ;
        RECT  0.575 1.180 1.050 1.285 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.310 1.330 0.940 ;
        RECT  0.750 0.310 1.240 0.400 ;
        RECT  0.650 0.310 0.750 0.890 ;
        RECT  0.480 0.780 0.650 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.165 1.600 0.165 ;
        RECT  1.420 -0.165 1.520 0.695 ;
        RECT  0.425 -0.165 1.420 0.165 ;
        RECT  0.425 0.300 0.525 0.400 ;
        RECT  0.315 -0.165 0.425 0.400 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.635 1.600 1.965 ;
        RECT  1.405 1.040 1.515 1.965 ;
        RECT  0.770 1.635 1.405 1.965 ;
        RECT  0.770 1.400 1.035 1.500 ;
        RECT  0.630 1.400 0.770 1.965 ;
        RECT  0.315 1.400 0.630 1.500 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.840 0.755 0.940 1.090 ;
        RECT  0.390 1.000 0.840 1.090 ;
        RECT  0.300 0.510 0.390 1.290 ;
        RECT  0.055 0.510 0.300 0.600 ;
        RECT  0.055 1.200 0.300 1.290 ;
    END
END IND2D2

MACRO IND2D4
    CLASS CORE ;
    FOREIGN IND2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.510 2.875 0.680 ;
        RECT  2.725 1.040 2.835 1.470 ;
        RECT  2.650 1.040 2.725 1.210 ;
        RECT  2.350 0.510 2.650 1.210 ;
        RECT  2.165 0.510 2.350 0.620 ;
        RECT  2.315 1.040 2.350 1.210 ;
        RECT  2.205 1.040 2.315 1.470 ;
        RECT  1.795 1.040 2.205 1.210 ;
        RECT  1.685 1.040 1.795 1.470 ;
        RECT  1.275 1.040 1.685 1.210 ;
        RECT  1.165 1.040 1.275 1.470 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 0.780 2.260 0.890 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.245 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.745 -0.165 3.200 0.165 ;
        RECT  1.745 0.310 1.845 0.420 ;
        RECT  1.635 -0.165 1.745 0.420 ;
        RECT  1.225 -0.165 1.635 0.165 ;
        RECT  1.225 0.310 1.325 0.420 ;
        RECT  1.115 -0.165 1.225 0.420 ;
        RECT  0.705 -0.165 1.115 0.165 ;
        RECT  0.595 -0.165 0.705 0.695 ;
        RECT  0.185 -0.165 0.595 0.165 ;
        RECT  0.075 -0.165 0.185 0.575 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.095 1.635 3.200 1.965 ;
        RECT  2.985 1.040 3.095 1.965 ;
        RECT  2.575 1.635 2.985 1.965 ;
        RECT  2.435 1.320 2.575 1.965 ;
        RECT  2.055 1.635 2.435 1.965 ;
        RECT  1.945 1.320 2.055 1.965 ;
        RECT  1.565 1.635 1.945 1.965 ;
        RECT  1.425 1.320 1.565 1.965 ;
        RECT  1.015 1.635 1.425 1.965 ;
        RECT  0.905 1.040 1.015 1.965 ;
        RECT  0.705 1.635 0.905 1.965 ;
        RECT  0.595 1.040 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.795 1.040 2.205 1.210 ;
        RECT  1.685 1.040 1.795 1.470 ;
        RECT  1.275 1.040 1.685 1.210 ;
        RECT  1.165 1.040 1.275 1.470 ;
        RECT  2.985 0.275 3.095 0.695 ;
        RECT  2.055 0.310 2.985 0.420 ;
        RECT  1.945 0.310 2.055 0.620 ;
        RECT  1.535 0.530 1.945 0.620 ;
        RECT  0.445 0.785 1.710 0.890 ;
        RECT  1.425 0.275 1.535 0.695 ;
        RECT  1.015 0.530 1.425 0.620 ;
        RECT  0.905 0.275 1.015 0.695 ;
        RECT  0.335 0.275 0.445 1.470 ;
        RECT  2.750 0.510 2.875 0.680 ;
        RECT  2.750 1.040 2.835 1.470 ;
        RECT  2.165 0.510 2.250 0.620 ;
        RECT  2.205 1.040 2.250 1.470 ;
    END
END IND2D4

MACRO IND3D0
    CLASS CORE ;
    FOREIGN IND3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1410 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.330 1.345 0.440 ;
        RECT  1.185 1.200 1.295 1.490 ;
        RECT  0.775 1.200 1.185 1.300 ;
        RECT  0.750 1.200 0.775 1.490 ;
        RECT  0.650 0.330 0.750 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.220 0.710 1.350 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.960 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.710 0.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.450 -0.165 1.400 0.165 ;
        RECT  0.450 0.310 0.550 0.420 ;
        RECT  0.340 -0.165 0.450 0.420 ;
        RECT  0.000 -0.165 0.340 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.985 1.635 1.400 1.965 ;
        RECT  0.985 1.390 1.085 1.500 ;
        RECT  0.875 1.390 0.985 1.965 ;
        RECT  0.450 1.635 0.875 1.965 ;
        RECT  0.450 1.380 0.550 1.490 ;
        RECT  0.340 1.380 0.450 1.965 ;
        RECT  0.000 1.635 0.340 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.460 0.530 0.560 1.270 ;
        RECT  0.225 0.530 0.460 0.620 ;
        RECT  0.225 1.180 0.460 1.270 ;
        RECT  0.115 0.275 0.225 0.620 ;
        RECT  0.115 1.180 0.225 1.490 ;
    END
END IND3D0

MACRO IND3D1
    CLASS CORE ;
    FOREIGN IND3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.490 1.345 0.600 ;
        RECT  0.775 1.200 1.345 1.300 ;
        RECT  0.750 1.200 0.775 1.400 ;
        RECT  0.650 0.490 0.750 1.400 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.090 ;
        RECT  1.210 0.710 1.250 0.940 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.960 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.210 0.710 0.250 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.450 -0.165 1.400 0.165 ;
        RECT  0.450 0.310 0.550 0.420 ;
        RECT  0.340 -0.165 0.450 0.420 ;
        RECT  0.000 -0.165 0.340 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.995 1.635 1.400 1.965 ;
        RECT  0.995 1.390 1.085 1.495 ;
        RECT  0.885 1.390 0.995 1.965 ;
        RECT  0.450 1.635 0.885 1.965 ;
        RECT  0.450 1.380 0.550 1.490 ;
        RECT  0.340 1.380 0.450 1.965 ;
        RECT  0.000 1.635 0.340 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.470 0.530 0.560 1.270 ;
        RECT  0.225 0.530 0.470 0.620 ;
        RECT  0.225 1.180 0.470 1.270 ;
        RECT  0.115 0.275 0.225 0.620 ;
        RECT  0.115 1.180 0.225 1.480 ;
    END
END IND3D1

MACRO IND3D2
    CLASS CORE ;
    FOREIGN IND3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.500 2.105 0.600 ;
        RECT  1.955 1.040 2.065 1.470 ;
        RECT  1.950 1.040 1.955 1.150 ;
        RECT  1.850 0.500 1.950 1.150 ;
        RECT  1.550 1.040 1.850 1.150 ;
        RECT  1.435 1.040 1.550 1.490 ;
        RECT  0.765 1.040 1.435 1.150 ;
        RECT  0.650 1.040 0.765 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.350 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.550 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.055 -0.165 2.400 0.165 ;
        RECT  0.945 -0.165 1.055 0.410 ;
        RECT  0.555 -0.165 0.945 0.165 ;
        RECT  0.865 0.305 0.945 0.410 ;
        RECT  0.445 -0.165 0.555 0.410 ;
        RECT  0.000 -0.165 0.445 0.165 ;
        RECT  0.345 0.305 0.445 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 1.635 2.400 1.965 ;
        RECT  2.215 1.040 2.325 1.965 ;
        RECT  1.805 1.635 2.215 1.965 ;
        RECT  1.695 1.260 1.805 1.965 ;
        RECT  1.285 1.635 1.695 1.965 ;
        RECT  1.175 1.260 1.285 1.965 ;
        RECT  1.025 1.635 1.175 1.965 ;
        RECT  0.915 1.260 1.025 1.965 ;
        RECT  0.505 1.635 0.915 1.965 ;
        RECT  0.395 1.260 0.505 1.965 ;
        RECT  0.000 1.635 0.395 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.215 0.305 2.325 0.585 ;
        RECT  1.145 0.305 2.215 0.410 ;
        RECT  0.620 0.520 1.595 0.620 ;
        RECT  0.530 0.780 0.815 0.890 ;
        RECT  0.440 0.500 0.530 1.150 ;
        RECT  0.085 0.500 0.440 0.600 ;
        RECT  0.245 1.040 0.440 1.150 ;
        RECT  0.135 1.040 0.245 1.470 ;
    END
END IND3D2

MACRO IND3D4
    CLASS CORE ;
    FOREIGN IND3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.500 3.905 0.600 ;
        RECT  3.745 1.040 3.855 1.470 ;
        RECT  3.450 1.040 3.745 1.150 ;
        RECT  3.350 0.500 3.450 1.150 ;
        RECT  3.225 0.500 3.350 1.490 ;
        RECT  3.150 0.500 3.225 1.150 ;
        RECT  2.815 1.040 3.150 1.150 ;
        RECT  2.705 1.040 2.815 1.470 ;
        RECT  2.295 1.040 2.705 1.150 ;
        RECT  2.185 1.040 2.295 1.470 ;
        RECT  1.495 1.040 2.185 1.150 ;
        RECT  1.385 1.040 1.495 1.470 ;
        RECT  0.975 1.040 1.385 1.150 ;
        RECT  0.850 1.040 0.975 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 0.770 4.045 0.900 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.770 2.845 0.900 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.770 0.240 0.900 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.570 -0.165 4.200 0.165 ;
        RECT  1.570 0.300 1.785 0.410 ;
        RECT  1.430 -0.165 1.570 0.410 ;
        RECT  0.715 -0.165 1.430 0.165 ;
        RECT  1.075 0.300 1.430 0.410 ;
        RECT  0.605 -0.165 0.715 0.695 ;
        RECT  0.195 -0.165 0.605 0.165 ;
        RECT  0.085 -0.165 0.195 0.585 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.115 1.635 4.200 1.965 ;
        RECT  4.005 1.040 4.115 1.965 ;
        RECT  3.595 1.635 4.005 1.965 ;
        RECT  3.485 1.260 3.595 1.965 ;
        RECT  3.075 1.635 3.485 1.965 ;
        RECT  2.965 1.260 3.075 1.965 ;
        RECT  2.565 1.635 2.965 1.965 ;
        RECT  2.435 1.260 2.565 1.965 ;
        RECT  2.035 1.635 2.435 1.965 ;
        RECT  1.925 1.260 2.035 1.965 ;
        RECT  1.755 1.635 1.925 1.965 ;
        RECT  1.635 1.260 1.755 1.965 ;
        RECT  1.235 1.635 1.635 1.965 ;
        RECT  1.125 1.260 1.235 1.965 ;
        RECT  0.715 1.635 1.125 1.965 ;
        RECT  0.605 1.040 0.715 1.965 ;
        RECT  0.195 1.635 0.605 1.965 ;
        RECT  0.085 1.260 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.550 0.500 3.905 0.600 ;
        RECT  3.745 1.040 3.855 1.470 ;
        RECT  3.550 1.040 3.745 1.150 ;
        RECT  2.815 1.040 3.050 1.150 ;
        RECT  2.705 1.040 2.815 1.470 ;
        RECT  2.295 1.040 2.705 1.150 ;
        RECT  2.185 1.040 2.295 1.470 ;
        RECT  1.495 1.040 2.185 1.150 ;
        RECT  1.385 1.040 1.495 1.470 ;
        RECT  0.975 1.040 1.385 1.150 ;
        RECT  0.850 1.040 0.975 1.490 ;
        RECT  1.895 0.305 4.155 0.410 ;
        RECT  0.825 0.500 2.865 0.600 ;
        RECT  0.455 0.785 1.555 0.890 ;
        RECT  0.345 0.275 0.455 1.470 ;
    END
END IND3D4

MACRO IND4D0
    CLASS CORE ;
    FOREIGN IND4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1380 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.310 1.550 0.490 ;
        RECT  1.265 0.310 1.340 1.120 ;
        RECT  1.250 0.310 1.265 1.490 ;
        RECT  1.155 1.030 1.250 1.490 ;
        RECT  0.750 1.030 1.155 1.120 ;
        RECT  0.635 1.030 0.750 1.490 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.710 1.550 1.090 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.160 0.920 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.510 0.950 0.920 ;
        RECT  0.810 0.730 0.850 0.920 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.180 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 -0.165 1.600 0.165 ;
        RECT  0.445 0.305 0.535 0.420 ;
        RECT  0.335 -0.165 0.445 0.420 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 1.635 1.600 1.965 ;
        RECT  1.415 1.280 1.525 1.965 ;
        RECT  1.005 1.635 1.415 1.965 ;
        RECT  0.895 1.280 1.005 1.965 ;
        RECT  0.535 1.635 0.895 1.965 ;
        RECT  0.425 1.390 0.535 1.965 ;
        RECT  0.335 1.390 0.425 1.495 ;
        RECT  0.000 1.635 0.425 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.360 0.780 0.620 0.890 ;
        RECT  0.270 0.510 0.360 1.300 ;
        RECT  0.225 0.510 0.270 0.600 ;
        RECT  0.225 1.210 0.270 1.300 ;
        RECT  0.115 0.275 0.225 0.600 ;
        RECT  0.115 1.210 0.225 1.480 ;
    END
END IND4D0

MACRO IND4D1
    CLASS CORE ;
    FOREIGN IND4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.310 1.550 0.490 ;
        RECT  1.250 0.310 1.340 1.120 ;
        RECT  0.585 1.030 1.250 1.120 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.565 0.920 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.510 0.950 0.920 ;
        RECT  0.810 0.730 0.850 0.920 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.160 0.920 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.180 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 -0.165 1.600 0.165 ;
        RECT  0.445 0.305 0.535 0.420 ;
        RECT  0.335 -0.165 0.445 0.420 ;
        RECT  0.000 -0.165 0.335 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.635 1.600 1.965 ;
        RECT  0.970 1.390 1.555 1.500 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.335 1.390 0.830 1.500 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.450 0.730 1.550 1.300 ;
        RECT  1.430 0.730 1.450 0.940 ;
        RECT  0.360 1.210 1.450 1.300 ;
        RECT  0.270 0.510 0.360 1.300 ;
        RECT  0.225 0.510 0.270 0.600 ;
        RECT  0.225 1.210 0.270 1.300 ;
        RECT  0.115 0.275 0.225 0.600 ;
        RECT  0.115 1.210 0.225 1.480 ;
    END
END IND4D1

MACRO IND4D2
    CLASS CORE ;
    FOREIGN IND4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.500 3.145 0.610 ;
        RECT  2.550 1.015 2.885 1.120 ;
        RECT  2.435 0.500 2.550 1.120 ;
        RECT  0.565 1.015 2.435 1.120 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.550 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.255 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.165 3.200 0.165 ;
        RECT  0.770 0.305 1.015 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.305 0.300 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.635 3.200 1.965 ;
        RECT  2.170 1.390 2.625 1.495 ;
        RECT  2.030 1.390 2.170 1.965 ;
        RECT  1.625 1.390 2.030 1.495 ;
        RECT  0.770 1.635 2.030 1.965 ;
        RECT  0.770 1.390 1.315 1.495 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.315 1.390 0.630 1.495 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.995 0.775 3.085 1.300 ;
        RECT  2.675 0.775 2.995 0.890 ;
        RECT  0.455 1.210 2.995 1.300 ;
        RECT  1.895 0.305 2.890 0.410 ;
        RECT  1.785 0.500 2.345 0.610 ;
        RECT  1.675 0.305 1.785 0.610 ;
        RECT  1.125 0.305 1.675 0.410 ;
        RECT  0.565 0.500 1.565 0.610 ;
        RECT  0.365 0.510 0.455 1.300 ;
        RECT  0.055 0.510 0.365 0.600 ;
        RECT  0.055 1.210 0.365 1.300 ;
    END
END IND4D2

MACRO IND4D4
    CLASS CORE ;
    FOREIGN IND4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.500 5.110 0.610 ;
        RECT  4.650 1.015 5.100 1.120 ;
        RECT  4.350 0.500 4.650 1.120 ;
        RECT  0.805 1.015 4.350 1.120 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.2198 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.770 1.555 0.900 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2185 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.770 2.750 0.900 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2185 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.770 3.750 0.900 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.680 0.190 0.940 ;
        RECT  0.050 0.680 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 -0.165 5.400 0.165 ;
        RECT  0.595 -0.165 0.705 0.695 ;
        RECT  0.185 -0.165 0.595 0.165 ;
        RECT  0.075 -0.165 0.185 0.560 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.635 5.400 1.965 ;
        RECT  4.570 1.390 5.340 1.500 ;
        RECT  4.430 1.390 4.570 1.965 ;
        RECT  3.860 1.390 4.430 1.500 ;
        RECT  3.370 1.635 4.430 1.965 ;
        RECT  3.370 1.390 3.550 1.500 ;
        RECT  3.230 1.390 3.370 1.965 ;
        RECT  2.820 1.390 3.230 1.500 ;
        RECT  2.170 1.635 3.230 1.965 ;
        RECT  2.170 1.390 2.510 1.500 ;
        RECT  2.030 1.390 2.170 1.965 ;
        RECT  1.685 1.390 2.030 1.500 ;
        RECT  0.970 1.635 2.030 1.965 ;
        RECT  0.970 1.390 1.285 1.500 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.545 1.390 0.830 1.500 ;
        RECT  0.185 1.635 0.830 1.965 ;
        RECT  0.075 1.210 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.750 0.500 5.110 0.610 ;
        RECT  4.750 1.015 5.100 1.120 ;
        RECT  0.805 1.015 4.250 1.120 ;
        RECT  5.210 0.305 5.320 0.585 ;
        RECT  5.220 0.775 5.310 1.300 ;
        RECT  4.770 0.775 5.220 0.890 ;
        RECT  0.445 1.210 5.220 1.300 ;
        RECT  3.080 0.305 5.210 0.410 ;
        RECT  1.780 0.500 4.070 0.600 ;
        RECT  1.465 0.305 2.770 0.410 ;
        RECT  1.355 0.305 1.465 0.680 ;
        RECT  0.805 0.305 1.355 0.410 ;
        RECT  0.335 0.275 0.445 1.300 ;
    END
END IND4D4

MACRO INR2D0
    CLASS CORE ;
    FOREIGN INR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0930 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.420 ;
        RECT  0.795 0.510 1.050 0.600 ;
        RECT  0.895 1.310 1.050 1.420 ;
        RECT  0.685 0.280 0.795 0.600 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.960 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.105 -0.165 1.200 0.165 ;
        RECT  0.995 -0.165 1.105 0.400 ;
        RECT  0.485 -0.165 0.995 0.165 ;
        RECT  0.895 0.290 0.995 0.400 ;
        RECT  0.485 0.310 0.585 0.420 ;
        RECT  0.375 -0.165 0.485 0.420 ;
        RECT  0.000 -0.165 0.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 1.635 1.200 1.965 ;
        RECT  0.485 1.380 0.585 1.490 ;
        RECT  0.375 1.380 0.485 1.965 ;
        RECT  0.000 1.635 0.375 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.575 0.750 0.680 0.920 ;
        RECT  0.485 0.530 0.575 1.270 ;
        RECT  0.275 0.530 0.485 0.620 ;
        RECT  0.275 1.180 0.485 1.270 ;
        RECT  0.165 0.280 0.275 0.620 ;
        RECT  0.165 1.180 0.275 1.490 ;
    END
END INR2D0

MACRO INR2D1
    CLASS CORE ;
    FOREIGN INR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.375 ;
        RECT  0.795 0.510 1.050 0.600 ;
        RECT  0.850 1.265 1.050 1.375 ;
        RECT  0.685 0.390 0.795 0.600 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.960 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.165 1.200 0.165 ;
        RECT  1.015 0.300 1.105 0.400 ;
        RECT  0.905 -0.165 1.015 0.400 ;
        RECT  0.485 -0.165 0.905 0.165 ;
        RECT  0.485 0.310 0.585 0.420 ;
        RECT  0.375 -0.165 0.485 0.420 ;
        RECT  0.000 -0.165 0.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.635 1.200 1.965 ;
        RECT  0.495 1.380 0.585 1.490 ;
        RECT  0.385 1.380 0.495 1.965 ;
        RECT  0.000 1.635 0.385 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.575 0.750 0.680 0.920 ;
        RECT  0.485 0.530 0.575 1.270 ;
        RECT  0.275 0.530 0.485 0.620 ;
        RECT  0.275 1.180 0.485 1.270 ;
        RECT  0.165 0.280 0.275 0.620 ;
        RECT  0.165 1.180 0.275 1.490 ;
    END
END INR2D1

MACRO INR2D2
    CLASS CORE ;
    FOREIGN INR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.510 1.305 0.620 ;
        RECT  1.050 0.510 1.150 1.290 ;
        RECT  0.575 0.510 1.050 0.600 ;
        RECT  0.840 1.200 1.050 1.290 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.710 0.955 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 -0.165 1.600 0.165 ;
        RECT  1.405 -0.165 1.515 0.585 ;
        RECT  0.770 -0.165 1.405 0.165 ;
        RECT  0.770 0.300 1.045 0.400 ;
        RECT  0.630 -0.165 0.770 0.400 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.315 0.300 0.630 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.635 1.600 1.965 ;
        RECT  1.420 1.035 1.520 1.965 ;
        RECT  0.425 1.635 1.420 1.965 ;
        RECT  0.425 1.400 0.525 1.500 ;
        RECT  0.315 1.400 0.425 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.730 1.330 1.490 ;
        RECT  0.730 1.400 1.240 1.490 ;
        RECT  0.640 0.775 0.730 1.490 ;
        RECT  0.465 0.775 0.640 0.890 ;
        RECT  0.375 0.510 0.465 1.290 ;
        RECT  0.055 0.510 0.375 0.600 ;
        RECT  0.055 1.200 0.375 1.290 ;
    END
END INR2D2

MACRO INR2D4
    CLASS CORE ;
    FOREIGN INR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.300 2.750 1.410 ;
        RECT  0.815 0.300 2.650 0.410 ;
        RECT  1.050 1.280 2.650 1.410 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 0.710 2.350 0.890 ;
        RECT  2.050 0.710 2.150 1.085 ;
        RECT  1.350 0.985 2.050 1.085 ;
        RECT  1.250 0.710 1.350 1.085 ;
        RECT  1.050 0.710 1.250 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.190 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 -0.165 2.800 0.165 ;
        RECT  0.595 -0.165 0.705 0.685 ;
        RECT  0.185 -0.165 0.595 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.635 2.800 1.965 ;
        RECT  0.595 1.105 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.450 0.500 2.560 0.920 ;
        RECT  1.760 0.500 2.450 0.600 ;
        RECT  1.580 0.500 1.760 0.895 ;
        RECT  0.950 0.500 1.580 0.600 ;
        RECT  0.850 0.500 0.950 0.885 ;
        RECT  0.445 0.785 0.850 0.885 ;
        RECT  0.335 0.275 0.445 1.470 ;
    END
END INR2D4

MACRO INR2XD0
    CLASS CORE ;
    FOREIGN INR2XD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.420 ;
        RECT  0.795 0.510 1.050 0.600 ;
        RECT  0.895 1.310 1.050 1.420 ;
        RECT  0.685 0.280 0.795 0.600 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.710 0.960 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.105 -0.165 1.200 0.165 ;
        RECT  0.995 -0.165 1.105 0.400 ;
        RECT  0.485 -0.165 0.995 0.165 ;
        RECT  0.895 0.290 0.995 0.400 ;
        RECT  0.485 0.310 0.585 0.420 ;
        RECT  0.375 -0.165 0.485 0.420 ;
        RECT  0.000 -0.165 0.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 1.635 1.200 1.965 ;
        RECT  0.485 1.380 0.585 1.490 ;
        RECT  0.375 1.380 0.485 1.965 ;
        RECT  0.000 1.635 0.375 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.575 0.750 0.680 0.920 ;
        RECT  0.485 0.530 0.575 1.270 ;
        RECT  0.275 0.530 0.485 0.620 ;
        RECT  0.275 1.180 0.485 1.270 ;
        RECT  0.165 0.280 0.275 0.620 ;
        RECT  0.165 1.180 0.275 1.490 ;
    END
END INR2XD0

MACRO INR2XD1
    CLASS CORE ;
    FOREIGN INR2XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.290 1.255 0.600 ;
        RECT  1.145 0.290 1.150 1.310 ;
        RECT  1.050 0.510 1.145 1.310 ;
        RECT  0.735 0.510 1.050 0.600 ;
        RECT  0.840 1.200 1.050 1.310 ;
        RECT  0.625 0.290 0.735 0.600 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.710 0.955 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 -0.165 1.600 0.165 ;
        RECT  1.405 -0.165 1.515 0.490 ;
        RECT  0.945 -0.165 1.405 0.165 ;
        RECT  0.945 0.310 1.045 0.420 ;
        RECT  0.835 -0.165 0.945 0.420 ;
        RECT  0.425 -0.165 0.835 0.165 ;
        RECT  0.425 0.305 0.525 0.415 ;
        RECT  0.315 -0.165 0.425 0.415 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.635 1.600 1.965 ;
        RECT  1.420 1.040 1.520 1.965 ;
        RECT  0.425 1.635 1.420 1.965 ;
        RECT  0.425 1.390 0.525 1.500 ;
        RECT  0.315 1.390 0.425 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.730 1.330 1.510 ;
        RECT  0.730 1.420 1.240 1.510 ;
        RECT  0.640 0.775 0.730 1.510 ;
        RECT  0.465 0.775 0.640 0.890 ;
        RECT  0.375 0.505 0.465 1.300 ;
        RECT  0.055 0.505 0.375 0.600 ;
        RECT  0.055 1.200 0.375 1.300 ;
    END
END INR2XD1

MACRO INR2XD2
    CLASS CORE ;
    FOREIGN INR2XD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 0.280 2.265 0.600 ;
        RECT  2.150 0.475 2.155 0.600 ;
        RECT  2.050 0.475 2.150 1.290 ;
        RECT  1.750 0.475 2.050 0.565 ;
        RECT  1.850 1.180 2.050 1.290 ;
        RECT  1.635 0.280 1.750 0.565 ;
        RECT  1.225 0.475 1.635 0.565 ;
        RECT  1.115 0.280 1.225 0.565 ;
        RECT  0.850 0.475 1.115 0.565 ;
        RECT  0.850 1.110 1.015 1.290 ;
        RECT  0.745 0.475 0.850 1.290 ;
        RECT  0.705 0.475 0.745 0.565 ;
        RECT  0.595 0.280 0.705 0.565 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.1716 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.675 1.950 0.890 ;
        RECT  1.055 0.675 1.650 0.765 ;
        RECT  0.945 0.675 1.055 0.940 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.525 -0.165 2.600 0.165 ;
        RECT  2.415 -0.165 2.525 0.490 ;
        RECT  1.955 -0.165 2.415 0.165 ;
        RECT  1.955 0.275 2.055 0.385 ;
        RECT  1.845 -0.165 1.955 0.385 ;
        RECT  1.435 -0.165 1.845 0.165 ;
        RECT  1.435 0.275 1.535 0.385 ;
        RECT  1.325 -0.165 1.435 0.385 ;
        RECT  0.915 -0.165 1.325 0.165 ;
        RECT  0.915 0.275 1.015 0.385 ;
        RECT  0.805 -0.165 0.915 0.385 ;
        RECT  0.395 -0.165 0.805 0.165 ;
        RECT  0.395 0.300 0.495 0.410 ;
        RECT  0.285 -0.165 0.395 0.410 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.525 1.635 2.600 1.965 ;
        RECT  2.425 1.060 2.525 1.965 ;
        RECT  1.485 1.635 2.425 1.965 ;
        RECT  1.375 1.310 1.485 1.965 ;
        RECT  0.475 1.635 1.375 1.965 ;
        RECT  0.365 1.380 0.475 1.965 ;
        RECT  0.285 1.380 0.365 1.490 ;
        RECT  0.000 1.635 0.365 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.330 0.750 2.380 0.920 ;
        RECT  2.240 0.750 2.330 1.490 ;
        RECT  1.735 1.400 2.240 1.490 ;
        RECT  1.625 1.090 1.735 1.490 ;
        RECT  1.535 1.090 1.625 1.200 ;
        RECT  1.325 0.855 1.535 1.200 ;
        RECT  1.245 1.090 1.325 1.200 ;
        RECT  1.135 1.090 1.245 1.490 ;
        RECT  0.655 1.400 1.135 1.490 ;
        RECT  0.565 0.780 0.655 1.490 ;
        RECT  0.435 0.780 0.565 0.890 ;
        RECT  0.345 0.510 0.435 1.290 ;
        RECT  0.185 0.510 0.345 0.600 ;
        RECT  0.185 1.200 0.345 1.290 ;
        RECT  0.075 0.355 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.390 ;
    END
END INR2XD2

MACRO INR2XD4
    CLASS CORE ;
    FOREIGN INR2XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.095 4.135 1.265 ;
        RECT  2.935 0.275 3.045 0.655 ;
        RECT  2.850 0.545 2.935 0.655 ;
        RECT  2.550 0.545 2.850 1.265 ;
        RECT  2.525 0.545 2.550 0.655 ;
        RECT  2.365 1.095 2.550 1.265 ;
        RECT  2.415 0.275 2.525 0.655 ;
        RECT  2.005 0.545 2.415 0.655 ;
        RECT  1.895 0.275 2.005 0.655 ;
        RECT  1.485 0.545 1.895 0.655 ;
        RECT  1.375 0.275 1.485 0.655 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.3432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.780 2.110 0.890 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.025 0.710 5.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.165 5.200 0.165 ;
        RECT  5.015 -0.165 5.125 0.585 ;
        RECT  4.605 -0.165 5.015 0.165 ;
        RECT  4.495 -0.165 4.605 0.670 ;
        RECT  3.305 -0.165 4.495 0.165 ;
        RECT  3.195 -0.165 3.305 0.670 ;
        RECT  2.785 -0.165 3.195 0.165 ;
        RECT  2.675 -0.165 2.785 0.455 ;
        RECT  2.265 -0.165 2.675 0.165 ;
        RECT  2.135 -0.165 2.265 0.455 ;
        RECT  1.765 -0.165 2.135 0.165 ;
        RECT  1.635 -0.165 1.765 0.455 ;
        RECT  1.225 -0.165 1.635 0.165 ;
        RECT  1.115 -0.165 1.225 0.670 ;
        RECT  0.000 -0.165 1.115 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.635 5.200 1.965 ;
        RECT  5.015 1.200 5.125 1.965 ;
        RECT  4.605 1.635 5.015 1.965 ;
        RECT  4.495 1.060 4.605 1.965 ;
        RECT  2.005 1.635 4.495 1.965 ;
        RECT  1.895 1.260 2.005 1.965 ;
        RECT  1.485 1.635 1.895 1.965 ;
        RECT  1.375 1.260 1.485 1.965 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.855 1.260 0.965 1.965 ;
        RECT  0.445 1.635 0.855 1.965 ;
        RECT  0.335 1.260 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 1.095 4.135 1.265 ;
        RECT  2.950 0.275 3.045 0.655 ;
        RECT  2.415 0.275 2.450 0.655 ;
        RECT  2.365 1.095 2.450 1.265 ;
        RECT  2.005 0.545 2.415 0.655 ;
        RECT  1.895 0.275 2.005 0.655 ;
        RECT  1.485 0.545 1.895 0.655 ;
        RECT  1.375 0.275 1.485 0.655 ;
        RECT  4.755 0.275 4.865 1.490 ;
        RECT  3.135 0.780 4.755 0.890 ;
        RECT  2.265 1.375 4.395 1.485 ;
        RECT  2.155 1.040 2.265 1.485 ;
        RECT  1.745 1.040 2.155 1.150 ;
        RECT  1.635 1.040 1.745 1.495 ;
        RECT  1.225 1.040 1.635 1.150 ;
        RECT  1.115 1.040 1.225 1.495 ;
        RECT  0.705 1.040 1.115 1.150 ;
        RECT  0.595 1.040 0.705 1.495 ;
        RECT  0.185 1.040 0.595 1.150 ;
        RECT  0.075 1.040 0.185 1.495 ;
    END
END INR2XD4

MACRO INR3D0
    CLASS CORE ;
    FOREIGN INR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1870 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.350 1.310 ;
        RECT  1.245 0.510 1.250 0.600 ;
        RECT  1.085 1.200 1.250 1.310 ;
        RECT  1.135 0.285 1.245 0.600 ;
        RECT  0.725 0.510 1.135 0.600 ;
        RECT  0.615 0.285 0.725 0.600 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.155 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 0.710 0.820 0.940 ;
        RECT  0.645 0.710 0.755 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 -0.165 1.400 0.165 ;
        RECT  0.935 0.310 1.035 0.420 ;
        RECT  0.825 -0.165 0.935 0.420 ;
        RECT  0.415 -0.165 0.825 0.165 ;
        RECT  0.415 0.310 0.515 0.420 ;
        RECT  0.305 -0.165 0.415 0.420 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.415 1.635 1.400 1.965 ;
        RECT  0.415 1.380 0.515 1.490 ;
        RECT  0.305 1.380 0.415 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.430 0.750 0.555 0.920 ;
        RECT  0.340 0.510 0.430 1.290 ;
        RECT  0.205 0.510 0.340 0.600 ;
        RECT  0.205 1.200 0.340 1.290 ;
        RECT  0.095 0.285 0.205 0.600 ;
        RECT  0.095 1.200 0.205 1.480 ;
    END
END INR3D0

MACRO INR3D1
    CLASS CORE ;
    FOREIGN INR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.520 1.105 0.620 ;
        RECT  0.150 1.190 1.025 1.290 ;
        RECT  0.050 0.520 0.150 1.290 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.310 1.365 0.690 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.800 1.370 0.890 ;
        RECT  0.850 0.710 1.150 0.890 ;
        RECT  0.470 0.775 0.850 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 1.950 1.090 ;
        RECT  1.680 0.780 1.850 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.705 -0.165 2.000 0.165 ;
        RECT  1.595 -0.165 1.705 0.415 ;
        RECT  0.570 -0.165 1.595 0.165 ;
        RECT  1.505 0.305 1.595 0.415 ;
        RECT  0.570 0.305 0.845 0.410 ;
        RECT  0.430 -0.165 0.570 0.410 ;
        RECT  0.000 -0.165 0.430 0.165 ;
        RECT  0.410 0.290 0.430 0.410 ;
        RECT  0.075 0.290 0.410 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.635 2.000 1.965 ;
        RECT  0.970 1.400 1.705 1.495 ;
        RECT  0.830 1.400 0.970 1.965 ;
        RECT  0.045 1.400 0.830 1.495 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.815 0.375 1.925 0.600 ;
        RECT  1.815 1.200 1.925 1.410 ;
        RECT  1.580 0.510 1.815 0.600 ;
        RECT  1.580 1.200 1.815 1.290 ;
        RECT  1.480 0.510 1.580 1.290 ;
        RECT  1.475 1.000 1.480 1.290 ;
        RECT  0.365 1.000 1.475 1.090 ;
        RECT  0.260 0.730 0.365 1.090 ;
    END
END INR3D1

MACRO INR3D2
    CLASS CORE ;
    FOREIGN INR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3380 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.505 2.150 1.490 ;
        RECT  1.750 0.505 2.050 0.605 ;
        RECT  1.105 1.390 2.050 1.490 ;
        RECT  0.765 0.510 1.750 0.600 ;
        RECT  0.650 0.310 0.765 0.600 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.710 1.630 0.920 ;
        RECT  1.450 0.710 1.545 1.085 ;
        RECT  0.950 0.995 1.450 1.085 ;
        RECT  0.855 0.710 0.950 1.085 ;
        RECT  0.760 0.710 0.855 0.920 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.780 0.290 0.890 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.095 -0.165 2.200 0.165 ;
        RECT  1.925 -0.165 2.095 0.405 ;
        RECT  1.575 -0.165 1.925 0.165 ;
        RECT  1.405 -0.165 1.575 0.405 ;
        RECT  1.055 -0.165 1.405 0.165 ;
        RECT  0.885 -0.165 1.055 0.405 ;
        RECT  0.535 -0.165 0.885 0.165 ;
        RECT  0.365 -0.165 0.535 0.405 ;
        RECT  0.000 -0.165 0.365 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.535 1.635 2.200 1.965 ;
        RECT  0.365 1.395 0.535 1.965 ;
        RECT  0.000 1.635 0.365 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.780 0.710 1.910 1.300 ;
        RECT  0.510 1.195 1.780 1.300 ;
        RECT  0.510 0.750 0.590 0.920 ;
        RECT  0.420 0.510 0.510 1.300 ;
        RECT  0.245 0.510 0.420 0.600 ;
        RECT  0.245 1.200 0.420 1.300 ;
        RECT  0.130 0.320 0.245 0.600 ;
        RECT  0.135 1.200 0.245 1.470 ;
    END
END INR3D2

MACRO INR3D4
    CLASS CORE ;
    FOREIGN INR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.285 3.750 1.505 ;
        RECT  0.785 0.285 3.650 0.390 ;
        RECT  1.285 1.360 3.650 1.505 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.660 2.960 1.090 ;
        RECT  2.380 0.660 2.850 0.750 ;
        RECT  2.290 0.660 2.380 1.090 ;
        RECT  2.020 1.000 2.290 1.090 ;
        RECT  1.930 0.660 2.020 1.090 ;
        RECT  1.550 0.660 1.930 0.750 ;
        RECT  1.440 0.660 1.550 1.090 ;
        RECT  1.295 0.750 1.440 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2203 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.220 0.710 3.350 1.270 ;
        RECT  2.640 1.180 3.220 1.270 ;
        RECT  2.470 0.840 2.640 1.270 ;
        RECT  1.840 1.180 2.470 1.270 ;
        RECT  1.650 0.840 1.840 1.270 ;
        RECT  1.150 1.180 1.650 1.270 ;
        RECT  1.050 0.710 1.150 1.270 ;
        RECT  0.990 0.710 1.050 0.920 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.190 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 3.800 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.635 3.800 1.965 ;
        RECT  0.075 1.220 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.450 0.480 3.560 0.920 ;
        RECT  2.200 0.480 3.450 0.570 ;
        RECT  2.110 0.480 2.200 0.890 ;
        RECT  0.810 0.480 2.110 0.570 ;
        RECT  0.665 0.480 0.810 0.905 ;
        RECT  0.445 0.765 0.665 0.905 ;
        RECT  0.335 0.275 0.445 1.470 ;
    END
END INR3D4

MACRO INR4D0
    CLASS CORE ;
    FOREIGN INR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1740 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.310 ;
        RECT  1.245 0.510 1.450 0.600 ;
        RECT  1.345 1.200 1.450 1.310 ;
        RECT  1.135 0.285 1.245 0.600 ;
        RECT  0.725 0.510 1.135 0.600 ;
        RECT  0.615 0.285 0.725 0.600 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.970 0.710 1.050 0.940 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.940 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.550 -0.165 1.600 0.165 ;
        RECT  1.440 -0.165 1.550 0.400 ;
        RECT  0.935 -0.165 1.440 0.165 ;
        RECT  1.345 0.290 1.440 0.400 ;
        RECT  0.935 0.310 1.035 0.420 ;
        RECT  0.825 -0.165 0.935 0.420 ;
        RECT  0.415 -0.165 0.825 0.165 ;
        RECT  0.415 0.310 0.515 0.420 ;
        RECT  0.305 -0.165 0.415 0.420 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.415 1.635 1.600 1.965 ;
        RECT  0.415 1.380 0.515 1.490 ;
        RECT  0.305 1.380 0.415 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.430 0.750 0.555 0.920 ;
        RECT  0.340 0.510 0.430 1.290 ;
        RECT  0.205 0.510 0.340 0.600 ;
        RECT  0.205 1.200 0.340 1.290 ;
        RECT  0.095 0.285 0.205 0.600 ;
        RECT  0.095 1.200 0.205 1.480 ;
    END
END INR4D0

MACRO INR4D1
    CLASS CORE ;
    FOREIGN INR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3270 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.500 2.555 0.600 ;
        RECT  1.550 1.015 2.125 1.115 ;
        RECT  1.450 0.500 1.550 1.115 ;
        RECT  0.595 0.500 1.450 0.610 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0763 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.165 0.890 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.400 0.710 2.550 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.300 -0.165 2.600 0.165 ;
        RECT  2.125 -0.165 2.300 0.410 ;
        RECT  0.770 -0.165 2.125 0.165 ;
        RECT  0.770 0.310 1.065 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.315 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.635 2.600 1.965 ;
        RECT  0.770 1.385 1.265 1.485 ;
        RECT  0.630 1.385 0.770 1.965 ;
        RECT  0.525 1.385 0.630 1.485 ;
        RECT  0.000 1.635 0.630 1.965 ;
        RECT  0.315 1.380 0.525 1.485 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.595 1.205 2.555 1.295 ;
        RECT  1.105 0.730 1.215 1.115 ;
        RECT  0.430 1.005 1.105 1.115 ;
        RECT  0.340 0.510 0.430 1.290 ;
        RECT  0.205 0.510 0.340 0.600 ;
        RECT  0.205 1.200 0.340 1.290 ;
        RECT  0.095 0.275 0.205 0.600 ;
        RECT  0.095 1.200 0.205 1.480 ;
    END
END INR4D1

MACRO INR4D2
    CLASS CORE ;
    FOREIGN INR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.425 3.960 1.490 ;
        RECT  0.820 0.425 3.850 0.525 ;
        RECT  3.280 1.380 3.850 1.490 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.640 3.750 0.890 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.640 2.960 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.640 2.160 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.220 0.890 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 -0.165 4.400 0.165 ;
        RECT  4.000 -0.165 4.170 0.335 ;
        RECT  3.575 -0.165 4.000 0.165 ;
        RECT  3.405 -0.165 3.575 0.335 ;
        RECT  3.005 -0.165 3.405 0.165 ;
        RECT  2.835 -0.165 3.005 0.335 ;
        RECT  2.435 -0.165 2.835 0.165 ;
        RECT  2.265 -0.165 2.435 0.335 ;
        RECT  1.865 -0.165 2.265 0.165 ;
        RECT  1.695 -0.165 1.865 0.335 ;
        RECT  1.295 -0.165 1.695 0.165 ;
        RECT  1.125 -0.165 1.295 0.335 ;
        RECT  0.720 -0.165 1.125 0.165 ;
        RECT  0.610 -0.165 0.720 0.520 ;
        RECT  0.185 -0.165 0.610 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.635 4.400 1.965 ;
        RECT  1.250 1.220 1.360 1.965 ;
        RECT  0.840 1.635 1.250 1.965 ;
        RECT  0.730 1.000 0.840 1.965 ;
        RECT  0.185 1.635 0.730 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.180 1.000 3.750 1.110 ;
        RECT  3.070 1.000 3.180 1.430 ;
        RECT  2.500 1.000 3.070 1.110 ;
        RECT  2.400 1.320 2.970 1.430 ;
        RECT  2.290 1.000 2.400 1.430 ;
        RECT  1.720 1.320 2.290 1.430 ;
        RECT  1.620 1.000 2.190 1.110 ;
        RECT  1.510 1.000 1.620 1.430 ;
        RECT  1.100 1.000 1.510 1.110 ;
        RECT  0.445 0.650 1.475 0.760 ;
        RECT  0.990 1.000 1.100 1.430 ;
        RECT  0.335 0.335 0.445 1.470 ;
    END
END INR4D2

MACRO INR4D4
    CLASS CORE ;
    FOREIGN INR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.500 5.115 0.620 ;
        RECT  4.850 1.040 5.115 1.210 ;
        RECT  4.550 0.500 4.850 1.210 ;
        RECT  1.025 0.500 4.550 0.620 ;
        RECT  4.385 1.040 4.550 1.210 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.2188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.960 0.710 5.350 0.920 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2198 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.710 4.000 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2186 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.710 2.740 0.890 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1098 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.710 0.220 0.890 ;
        RECT  0.050 0.710 0.155 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.970 -0.165 5.400 0.165 ;
        RECT  4.970 0.300 5.355 0.410 ;
        RECT  4.830 -0.165 4.970 0.410 ;
        RECT  3.770 -0.165 4.830 0.165 ;
        RECT  4.645 0.300 4.830 0.410 ;
        RECT  3.770 0.305 4.340 0.410 ;
        RECT  3.630 -0.165 3.770 0.410 ;
        RECT  2.170 -0.165 3.630 0.165 ;
        RECT  2.905 0.305 3.630 0.410 ;
        RECT  2.170 0.300 2.515 0.410 ;
        RECT  2.030 -0.165 2.170 0.410 ;
        RECT  0.925 -0.165 2.030 0.165 ;
        RECT  1.785 0.300 2.030 0.410 ;
        RECT  0.815 -0.165 0.925 0.675 ;
        RECT  0.705 -0.165 0.815 0.165 ;
        RECT  0.595 -0.165 0.705 0.675 ;
        RECT  0.185 -0.165 0.595 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.185 1.635 5.400 1.965 ;
        RECT  1.075 1.260 1.185 1.965 ;
        RECT  0.185 1.635 1.075 1.965 ;
        RECT  0.075 1.260 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.950 0.500 5.115 0.620 ;
        RECT  4.950 1.040 5.115 1.210 ;
        RECT  1.025 0.500 4.450 0.620 ;
        RECT  4.385 1.040 4.450 1.210 ;
        RECT  4.285 1.355 5.355 1.465 ;
        RECT  4.175 1.050 4.285 1.465 ;
        RECT  3.105 1.355 4.175 1.465 ;
        RECT  2.045 1.090 4.075 1.200 ;
        RECT  1.945 1.355 3.015 1.465 ;
        RECT  1.835 1.040 1.945 1.500 ;
        RECT  1.445 1.040 1.835 1.150 ;
        RECT  0.445 0.780 1.720 0.890 ;
        RECT  1.335 1.040 1.445 1.500 ;
        RECT  0.925 1.040 1.335 1.150 ;
        RECT  0.815 1.040 0.925 1.500 ;
        RECT  0.335 0.275 0.445 1.500 ;
    END
END INR4D4

MACRO INVD0
    CLASS CORE ;
    FOREIGN INVD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.440 0.550 1.360 ;
        RECT  0.295 0.440 0.440 0.550 ;
        RECT  0.295 1.250 0.440 1.360 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.705 0.350 1.095 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.165 0.600 0.165 ;
        RECT  0.085 -0.165 0.195 0.595 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 1.635 0.600 1.965 ;
        RECT  0.085 1.200 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END INVD0

MACRO INVD1
    CLASS CORE ;
    FOREIGN INVD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.275 0.550 1.490 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.190 1.120 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.250 -0.165 0.600 0.165 ;
        RECT  0.140 -0.165 0.250 0.560 ;
        RECT  0.000 -0.165 0.140 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.250 1.635 0.600 1.965 ;
        RECT  0.140 1.240 0.250 1.965 ;
        RECT  0.000 1.635 0.140 1.965 ;
        END
    END VDD
END INVD1

MACRO INVD12
    CLASS CORE ;
    FOREIGN INVD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.0920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.325 3.115 0.690 ;
        RECT  2.050 1.100 3.115 1.475 ;
        RECT  1.550 0.325 2.050 1.475 ;
        RECT  0.325 0.325 1.550 0.690 ;
        RECT  0.355 1.100 1.550 1.475 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.6618 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.800 1.340 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 -0.165 3.400 0.165 ;
        RECT  3.215 -0.165 3.330 0.690 ;
        RECT  0.215 -0.165 3.215 0.165 ;
        RECT  0.085 -0.165 0.215 0.595 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 1.635 3.400 1.965 ;
        RECT  3.215 1.080 3.330 1.965 ;
        RECT  0.215 1.635 3.215 1.965 ;
        RECT  0.085 1.200 0.215 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.150 0.325 3.115 0.690 ;
        RECT  2.150 1.100 3.115 1.475 ;
        RECT  0.325 0.325 1.450 0.690 ;
        RECT  0.355 1.100 1.450 1.475 ;
        RECT  2.210 0.800 3.170 0.940 ;
    END
END INVD12

MACRO INVD16
    CLASS CORE ;
    FOREIGN INVD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.4560 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.325 4.115 0.690 ;
        RECT  2.450 1.100 4.115 1.475 ;
        RECT  1.950 0.325 2.450 1.475 ;
        RECT  0.305 0.325 1.950 0.690 ;
        RECT  0.305 1.100 1.950 1.475 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.8828 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.800 1.790 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.690 ;
        RECT  0.185 -0.165 4.215 0.165 ;
        RECT  0.075 -0.165 0.185 0.595 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.055 4.325 1.965 ;
        RECT  0.185 1.635 4.215 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.325 4.115 0.690 ;
        RECT  2.550 1.100 4.115 1.475 ;
        RECT  0.305 0.325 1.850 0.690 ;
        RECT  0.305 1.100 1.850 1.475 ;
        RECT  2.640 0.800 4.170 0.940 ;
    END
END INVD16

MACRO INVD2
    CLASS CORE ;
    FOREIGN INVD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.605 0.550 1.130 ;
        RECT  0.425 0.275 0.455 1.470 ;
        RECT  0.345 0.275 0.425 0.695 ;
        RECT  0.345 1.040 0.425 1.470 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.165 0.800 0.165 ;
        RECT  0.605 -0.165 0.715 0.495 ;
        RECT  0.195 -0.165 0.605 0.165 ;
        RECT  0.085 -0.165 0.195 0.595 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.240 0.715 1.965 ;
        RECT  0.195 1.635 0.605 1.965 ;
        RECT  0.085 1.200 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END INVD2

MACRO INVD20
    CLASS CORE ;
    FOREIGN INVD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.8200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.325 5.095 0.690 ;
        RECT  2.850 1.100 5.095 1.475 ;
        RECT  2.350 0.325 2.850 1.475 ;
        RECT  0.305 0.325 2.350 0.690 ;
        RECT  0.305 1.100 2.350 1.475 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.1040 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.800 2.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.325 -0.165 5.400 0.165 ;
        RECT  5.215 -0.165 5.325 0.695 ;
        RECT  0.185 -0.165 5.215 0.165 ;
        RECT  0.075 -0.165 0.185 0.595 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.325 1.635 5.400 1.965 ;
        RECT  5.215 1.040 5.325 1.965 ;
        RECT  0.185 1.635 5.215 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.325 5.095 0.690 ;
        RECT  2.950 1.100 5.095 1.475 ;
        RECT  0.305 0.325 2.250 0.690 ;
        RECT  0.305 1.100 2.250 1.475 ;
        RECT  3.010 0.800 5.170 0.940 ;
    END
END INVD20

MACRO INVD24
    CLASS CORE ;
    FOREIGN INVD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 2.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.325 6.095 0.690 ;
        RECT  3.450 1.100 6.095 1.475 ;
        RECT  2.950 0.325 3.450 1.475 ;
        RECT  0.305 0.325 2.950 0.690 ;
        RECT  0.305 1.100 2.950 1.475 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.3250 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.800 2.790 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.325 -0.165 6.400 0.165 ;
        RECT  6.215 -0.165 6.325 0.695 ;
        RECT  0.185 -0.165 6.215 0.165 ;
        RECT  0.075 -0.165 0.185 0.595 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.325 1.635 6.400 1.965 ;
        RECT  6.215 1.040 6.325 1.965 ;
        RECT  0.185 1.635 6.215 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.550 0.325 6.095 0.690 ;
        RECT  3.550 1.100 6.095 1.475 ;
        RECT  0.305 0.325 2.850 0.690 ;
        RECT  0.305 1.100 2.850 1.475 ;
        RECT  3.610 0.800 6.040 0.940 ;
    END
END INVD24

MACRO INVD3
    CLASS CORE ;
    FOREIGN INVD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3690 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 0.275 1.045 1.470 ;
        RECT  0.550 0.650 0.920 0.950 ;
        RECT  0.415 0.275 0.550 1.490 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.785 -0.165 1.200 0.165 ;
        RECT  0.675 -0.165 0.785 0.540 ;
        RECT  0.265 -0.165 0.675 0.165 ;
        RECT  0.155 -0.165 0.265 0.595 ;
        RECT  0.000 -0.165 0.155 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.785 1.635 1.200 1.965 ;
        RECT  0.675 1.065 0.785 1.965 ;
        RECT  0.265 1.635 0.675 1.965 ;
        RECT  0.155 1.200 0.265 1.965 ;
        RECT  0.000 1.635 0.155 1.965 ;
        END
    END VDD
END INVD3

MACRO INVD4
    CLASS CORE ;
    FOREIGN INVD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.935 0.275 1.045 0.695 ;
        RECT  0.935 1.040 1.045 1.470 ;
        RECT  0.850 0.535 0.935 0.695 ;
        RECT  0.850 1.040 0.935 1.210 ;
        RECT  0.550 0.535 0.850 1.210 ;
        RECT  0.415 0.275 0.550 0.695 ;
        RECT  0.415 1.040 0.550 1.490 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.190 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 -0.165 1.400 0.165 ;
        RECT  1.195 -0.165 1.305 0.695 ;
        RECT  0.785 -0.165 1.195 0.165 ;
        RECT  0.675 -0.165 0.785 0.445 ;
        RECT  0.265 -0.165 0.675 0.165 ;
        RECT  0.155 -0.165 0.265 0.595 ;
        RECT  0.000 -0.165 0.155 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 1.635 1.400 1.965 ;
        RECT  1.195 1.040 1.305 1.965 ;
        RECT  0.785 1.635 1.195 1.965 ;
        RECT  0.675 1.300 0.785 1.965 ;
        RECT  0.265 1.635 0.675 1.965 ;
        RECT  0.155 1.200 0.265 1.965 ;
        RECT  0.000 1.635 0.155 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.275 1.045 0.695 ;
        RECT  0.950 1.040 1.045 1.470 ;
        RECT  0.415 0.275 0.450 0.695 ;
        RECT  0.415 1.040 0.450 1.490 ;
    END
END INVD4

MACRO INVD6
    CLASS CORE ;
    FOREIGN INVD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.275 1.475 0.695 ;
        RECT  1.340 1.040 1.475 1.490 ;
        RECT  1.050 0.525 1.340 0.695 ;
        RECT  1.050 1.040 1.340 1.210 ;
        RECT  0.965 0.525 1.050 1.210 ;
        RECT  0.835 0.275 0.965 1.490 ;
        RECT  0.750 0.525 0.835 1.210 ;
        RECT  0.455 0.525 0.750 0.695 ;
        RECT  0.455 1.040 0.750 1.210 ;
        RECT  0.325 0.275 0.455 0.695 ;
        RECT  0.325 1.040 0.455 1.490 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.3302 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.785 0.630 0.890 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.695 ;
        RECT  0.185 -0.165 1.615 0.165 ;
        RECT  0.075 -0.165 0.185 0.595 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.040 1.725 1.965 ;
        RECT  0.185 1.635 1.615 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.340 0.275 1.475 0.695 ;
        RECT  1.340 1.040 1.475 1.490 ;
        RECT  1.150 0.525 1.340 0.695 ;
        RECT  1.150 1.040 1.340 1.210 ;
        RECT  0.455 0.525 0.650 0.695 ;
        RECT  0.455 1.040 0.650 1.210 ;
        RECT  0.325 0.275 0.455 0.695 ;
        RECT  0.325 1.040 0.455 1.490 ;
    END
END INVD6

MACRO INVD8
    CLASS CORE ;
    FOREIGN INVD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.325 2.065 0.635 ;
        RECT  1.650 1.060 2.035 1.450 ;
        RECT  1.150 0.325 1.650 1.450 ;
        RECT  0.335 0.325 1.150 0.635 ;
        RECT  0.335 1.060 1.150 1.450 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.4368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.785 0.910 0.890 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 -0.165 2.400 0.165 ;
        RECT  2.185 -0.165 2.295 0.695 ;
        RECT  0.215 -0.165 2.185 0.165 ;
        RECT  0.105 -0.165 0.215 0.595 ;
        RECT  0.000 -0.165 0.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 1.635 2.400 1.965 ;
        RECT  2.185 1.040 2.295 1.965 ;
        RECT  0.215 1.635 2.185 1.965 ;
        RECT  0.105 1.200 0.215 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.750 0.325 2.065 0.635 ;
        RECT  1.750 1.060 2.035 1.450 ;
        RECT  0.335 0.325 1.050 0.635 ;
        RECT  0.335 1.060 1.050 1.450 ;
        RECT  1.760 0.785 2.140 0.900 ;
    END
END INVD8

MACRO IOA21D0
    CLASS CORE ;
    FOREIGN IOA21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0910 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.310 1.350 1.290 ;
        RECT  1.065 0.310 1.250 0.420 ;
        RECT  0.965 1.200 1.250 1.290 ;
        RECT  0.855 1.200 0.965 1.490 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.710 1.150 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.165 1.400 0.165 ;
        RECT  0.560 -0.165 0.740 0.405 ;
        RECT  0.000 -0.165 0.560 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.635 1.400 1.965 ;
        RECT  1.110 1.400 1.280 1.965 ;
        RECT  0.740 1.635 1.110 1.965 ;
        RECT  0.560 1.395 0.740 1.965 ;
        RECT  0.185 1.635 0.560 1.965 ;
        RECT  0.075 1.280 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.730 0.750 0.790 0.920 ;
        RECT  0.640 0.495 0.730 1.305 ;
        RECT  0.185 0.495 0.640 0.590 ;
        RECT  0.445 1.215 0.640 1.305 ;
        RECT  0.335 1.215 0.445 1.490 ;
        RECT  0.075 0.275 0.185 0.590 ;
    END
END IOA21D0

MACRO IOA21D1
    CLASS CORE ;
    FOREIGN IOA21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 0.490 1.350 1.300 ;
        RECT  1.250 0.400 1.290 1.300 ;
        RECT  1.180 0.400 1.250 0.590 ;
        RECT  1.005 1.210 1.250 1.300 ;
        RECT  0.895 1.210 1.005 1.480 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.700 1.150 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.565 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.210 0.940 ;
        RECT  0.050 0.700 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.775 -0.165 1.400 0.165 ;
        RECT  0.605 -0.165 0.775 0.405 ;
        RECT  0.000 -0.165 0.605 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.635 1.400 1.965 ;
        RECT  1.180 1.410 1.290 1.965 ;
        RECT  0.775 1.635 1.180 1.965 ;
        RECT  0.585 1.395 0.775 1.965 ;
        RECT  0.205 1.635 0.585 1.965 ;
        RECT  0.095 1.290 0.205 1.965 ;
        RECT  0.000 1.635 0.095 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.775 0.750 0.845 0.920 ;
        RECT  0.675 0.495 0.775 1.305 ;
        RECT  0.205 0.495 0.675 0.590 ;
        RECT  0.465 1.215 0.675 1.305 ;
        RECT  0.355 1.215 0.465 1.480 ;
        RECT  0.095 0.285 0.205 0.590 ;
    END
END IOA21D1

MACRO IOA21D2
    CLASS CORE ;
    FOREIGN IOA21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.355 1.075 1.465 1.485 ;
        RECT  1.350 1.075 1.355 1.305 ;
        RECT  1.250 0.485 1.350 1.305 ;
        RECT  1.080 0.485 1.250 0.590 ;
        RECT  0.965 1.215 1.250 1.305 ;
        RECT  0.865 1.215 0.965 1.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.700 1.150 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.565 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.210 0.940 ;
        RECT  0.050 0.700 0.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.755 -0.165 1.800 0.165 ;
        RECT  0.570 -0.165 0.755 0.405 ;
        RECT  0.000 -0.165 0.570 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.065 1.725 1.965 ;
        RECT  0.190 1.635 1.615 1.965 ;
        RECT  0.080 1.200 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.560 0.305 1.670 0.940 ;
        RECT  0.970 0.305 1.560 0.395 ;
        RECT  0.880 0.305 0.970 0.590 ;
        RECT  0.775 0.495 0.880 0.590 ;
        RECT  0.775 0.750 0.875 0.920 ;
        RECT  0.685 0.495 0.775 1.320 ;
        RECT  0.205 0.495 0.685 0.590 ;
        RECT  0.305 1.210 0.685 1.320 ;
        RECT  0.095 0.380 0.205 0.590 ;
    END
END IOA21D2

MACRO IOA21D4
    CLASS CORE ;
    FOREIGN IOA21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.695 1.460 ;
        RECT  2.350 0.495 2.555 1.210 ;
        RECT  1.995 0.495 2.350 0.660 ;
        RECT  2.145 1.040 2.350 1.210 ;
        RECT  2.035 1.040 2.145 1.460 ;
        RECT  0.945 1.205 2.035 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2194 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.550 0.890 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.710 0.950 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.245 0.930 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.660 -0.165 3.000 0.165 ;
        RECT  1.480 -0.165 1.660 0.410 ;
        RECT  0.000 -0.165 1.480 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.925 1.635 3.000 1.965 ;
        RECT  2.815 1.050 2.925 1.965 ;
        RECT  2.405 1.635 2.815 1.965 ;
        RECT  2.295 1.300 2.405 1.965 ;
        RECT  1.570 1.635 2.295 1.965 ;
        RECT  1.570 1.390 1.925 1.495 ;
        RECT  1.430 1.390 1.570 1.965 ;
        RECT  1.205 1.390 1.430 1.495 ;
        RECT  0.795 1.635 1.430 1.965 ;
        RECT  0.650 1.225 0.795 1.965 ;
        RECT  0.185 1.635 0.650 1.965 ;
        RECT  0.075 1.250 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.995 0.495 2.250 0.660 ;
        RECT  2.145 1.040 2.250 1.210 ;
        RECT  2.035 1.040 2.145 1.460 ;
        RECT  0.945 1.205 2.035 1.300 ;
        RECT  2.815 0.305 2.925 0.575 ;
        RECT  1.885 0.305 2.815 0.405 ;
        RECT  1.880 0.780 2.170 0.890 ;
        RECT  1.775 0.305 1.885 0.600 ;
        RECT  1.790 0.780 1.880 1.115 ;
        RECT  0.445 1.025 1.790 1.115 ;
        RECT  0.690 0.500 1.775 0.600 ;
        RECT  0.435 1.025 0.445 1.465 ;
        RECT  0.335 0.485 0.435 1.465 ;
        RECT  0.185 0.485 0.335 0.575 ;
        RECT  0.075 0.345 0.185 0.575 ;
    END
END IOA21D4

MACRO IOA22D0
    CLASS CORE ;
    FOREIGN IOA22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1190 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.210 1.750 1.490 ;
        RECT  0.980 1.210 1.615 1.300 ;
        RECT  0.965 0.285 0.980 1.300 ;
        RECT  0.880 0.285 0.965 1.490 ;
        RECT  0.835 0.285 0.880 0.490 ;
        RECT  0.850 1.110 0.880 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.710 1.640 0.940 ;
        RECT  1.450 0.710 1.550 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.180 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.165 1.800 0.165 ;
        RECT  1.320 -0.165 1.500 0.420 ;
        RECT  0.720 -0.165 1.320 0.165 ;
        RECT  0.540 -0.165 0.720 0.420 ;
        RECT  0.000 -0.165 0.540 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.635 1.800 1.965 ;
        RECT  1.080 1.390 1.260 1.965 ;
        RECT  0.740 1.635 1.080 1.965 ;
        RECT  0.560 1.380 0.740 1.965 ;
        RECT  0.185 1.635 0.560 1.965 ;
        RECT  0.075 1.290 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.615 0.285 1.725 0.600 ;
        RECT  1.205 0.510 1.615 0.600 ;
        RECT  1.095 0.285 1.205 0.600 ;
        RECT  0.730 0.750 0.790 0.920 ;
        RECT  0.640 0.510 0.730 1.290 ;
        RECT  0.185 0.510 0.640 0.600 ;
        RECT  0.445 1.200 0.640 1.290 ;
        RECT  0.335 1.200 0.445 1.480 ;
        RECT  0.075 0.290 0.185 0.600 ;
    END
END IOA22D0

MACRO IOA22D1
    CLASS CORE ;
    FOREIGN IOA22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2370 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.210 1.750 1.505 ;
        RECT  0.980 1.210 1.615 1.300 ;
        RECT  0.965 0.310 0.980 1.300 ;
        RECT  0.880 0.310 0.965 1.500 ;
        RECT  0.835 0.310 0.880 0.500 ;
        RECT  0.850 1.100 0.880 1.500 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.640 0.930 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.350 1.100 ;
        RECT  1.210 0.700 1.250 0.930 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.270 0.930 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.700 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.495 -0.165 1.800 0.165 ;
        RECT  1.325 -0.165 1.495 0.410 ;
        RECT  0.715 -0.165 1.325 0.165 ;
        RECT  0.545 -0.165 0.715 0.405 ;
        RECT  0.000 -0.165 0.545 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.255 1.635 1.800 1.965 ;
        RECT  1.085 1.390 1.255 1.965 ;
        RECT  0.735 1.635 1.085 1.965 ;
        RECT  0.565 1.395 0.735 1.965 ;
        RECT  0.185 1.635 0.565 1.965 ;
        RECT  0.075 1.290 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.615 0.370 1.725 0.590 ;
        RECT  1.205 0.500 1.615 0.590 ;
        RECT  1.095 0.370 1.205 0.590 ;
        RECT  0.730 0.750 0.790 0.920 ;
        RECT  0.640 0.500 0.730 1.305 ;
        RECT  0.185 0.500 0.640 0.590 ;
        RECT  0.445 1.215 0.640 1.305 ;
        RECT  0.335 1.215 0.445 1.480 ;
        RECT  0.075 0.290 0.185 0.590 ;
    END
END IOA22D1

MACRO IOA22D2
    CLASS CORE ;
    FOREIGN IOA22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.405 1.550 1.160 ;
        RECT  1.165 0.405 1.450 0.515 ;
        RECT  1.260 1.050 1.450 1.160 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.710 1.755 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0434 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.150 1.090 ;
        RECT  2.025 0.710 2.050 0.920 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.160 0.710 0.250 0.940 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.165 2.200 0.165 ;
        RECT  0.905 -0.165 1.015 0.515 ;
        RECT  0.185 -0.165 0.905 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.200 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 1.210 2.120 1.420 ;
        RECT  1.935 1.210 2.010 1.340 ;
        RECT  1.845 0.405 1.935 1.340 ;
        RECT  1.700 0.405 1.845 0.515 ;
        RECT  1.135 1.250 1.845 1.340 ;
        RECT  1.225 0.625 1.335 0.940 ;
        RECT  0.755 0.625 1.225 0.715 ;
        RECT  1.045 0.825 1.135 1.340 ;
        RECT  0.820 0.825 1.045 0.925 ;
        RECT  0.835 1.035 0.945 1.475 ;
        RECT  0.730 1.035 0.835 1.125 ;
        RECT  0.730 0.425 0.755 0.715 ;
        RECT  0.185 1.235 0.735 1.345 ;
        RECT  0.640 0.425 0.730 1.125 ;
        RECT  0.545 0.425 0.640 0.535 ;
        RECT  0.075 1.235 0.185 1.445 ;
    END
END IOA22D2

MACRO IOA22D4
    CLASS CORE ;
    FOREIGN IOA22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.015 2.795 1.125 ;
        RECT  2.650 0.310 2.750 0.635 ;
        RECT  2.635 0.310 2.650 1.125 ;
        RECT  2.350 0.525 2.635 1.125 ;
        RECT  2.065 0.525 2.350 0.635 ;
        RECT  2.065 1.015 2.350 1.125 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.150 1.090 ;
        RECT  2.990 0.710 3.050 0.940 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 3.550 1.090 ;
        RECT  3.420 0.710 3.450 0.940 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 1.150 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 -0.165 3.600 0.165 ;
        RECT  3.420 -0.165 3.525 0.485 ;
        RECT  3.005 -0.165 3.420 0.165 ;
        RECT  2.895 -0.165 3.005 0.490 ;
        RECT  2.170 -0.165 2.895 0.165 ;
        RECT  2.170 0.305 2.535 0.410 ;
        RECT  2.030 -0.165 2.170 0.410 ;
        RECT  0.485 -0.165 2.030 0.165 ;
        RECT  1.805 0.305 2.030 0.410 ;
        RECT  0.295 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.770 1.635 3.600 1.965 ;
        RECT  2.770 1.395 3.055 1.495 ;
        RECT  2.630 1.395 2.770 1.965 ;
        RECT  2.325 1.395 2.630 1.495 ;
        RECT  0.965 1.635 2.630 1.965 ;
        RECT  0.855 1.245 0.965 1.965 ;
        RECT  0.445 1.635 0.855 1.965 ;
        RECT  0.335 1.245 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 1.015 2.795 1.125 ;
        RECT  2.065 0.525 2.250 0.635 ;
        RECT  2.065 1.015 2.250 1.125 ;
        RECT  3.415 1.210 3.525 1.420 ;
        RECT  3.330 1.210 3.415 1.305 ;
        RECT  3.240 0.325 3.330 1.305 ;
        RECT  3.105 0.325 3.240 0.435 ;
        RECT  1.955 1.215 3.240 1.305 ;
        RECT  1.905 0.780 2.220 0.890 ;
        RECT  1.865 1.025 1.955 1.305 ;
        RECT  1.815 0.500 1.905 0.890 ;
        RECT  1.705 1.025 1.865 1.135 ;
        RECT  1.485 0.500 1.815 0.610 ;
        RECT  1.225 1.365 1.775 1.475 ;
        RECT  1.595 0.730 1.705 1.135 ;
        RECT  1.375 0.500 1.485 1.275 ;
        RECT  0.815 0.500 1.375 0.590 ;
        RECT  0.705 0.305 1.275 0.410 ;
        RECT  1.115 1.045 1.225 1.475 ;
        RECT  0.705 1.045 1.115 1.135 ;
        RECT  0.595 0.305 0.705 0.590 ;
        RECT  0.595 1.045 0.705 1.475 ;
        RECT  0.185 0.500 0.595 0.590 ;
        RECT  0.185 1.045 0.595 1.135 ;
        RECT  0.075 0.365 0.185 0.590 ;
        RECT  0.075 1.045 0.185 1.475 ;
    END
END IOA22D4

MACRO ISOHID1
    CLASS CORE ;
    FOREIGN ISOHID1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.300 1.150 1.500 ;
        RECT  0.995 0.300 1.050 0.685 ;
        RECT  0.995 1.100 1.050 1.500 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.780 0.660 0.890 ;
        RECT  0.450 0.710 0.550 1.100 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.755 0.350 0.920 ;
        RECT  0.050 0.500 0.150 0.920 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 -0.165 1.200 0.165 ;
        RECT  0.680 -0.165 0.850 0.390 ;
        RECT  0.270 -0.165 0.680 0.165 ;
        RECT  0.100 -0.165 0.270 0.390 ;
        RECT  0.000 -0.165 0.100 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.635 1.200 1.965 ;
        RECT  0.660 1.410 0.830 1.965 ;
        RECT  0.000 1.635 0.660 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 0.780 0.940 0.890 ;
        RECT  0.770 0.500 0.860 1.320 ;
        RECT  0.370 0.500 0.770 0.600 ;
        RECT  0.245 1.210 0.770 1.320 ;
        RECT  0.135 1.040 0.245 1.470 ;
    END
END ISOHID1

MACRO ISOHID2
    CLASS CORE ;
    FOREIGN ISOHID2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.575 1.150 1.170 ;
        RECT  0.940 0.295 1.050 0.685 ;
        RECT  1.040 1.060 1.050 1.170 ;
        RECT  0.930 1.060 1.040 1.470 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.605 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.240 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 -0.165 1.400 0.165 ;
        RECT  1.195 -0.165 1.315 0.475 ;
        RECT  0.795 -0.165 1.195 0.165 ;
        RECT  0.625 -0.165 0.795 0.390 ;
        RECT  0.210 -0.165 0.625 0.165 ;
        RECT  0.100 -0.165 0.210 0.590 ;
        RECT  0.000 -0.165 0.100 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 1.635 1.400 1.965 ;
        RECT  1.195 1.325 1.315 1.965 ;
        RECT  0.775 1.635 1.195 1.965 ;
        RECT  0.605 1.410 0.775 1.965 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.840 0.750 0.875 0.920 ;
        RECT  0.730 0.500 0.840 1.320 ;
        RECT  0.320 0.500 0.730 0.610 ;
        RECT  0.190 1.210 0.730 1.320 ;
        RECT  0.080 1.210 0.190 1.485 ;
    END
END ISOHID2

MACRO ISOHID4
    CLASS CORE ;
    FOREIGN ISOHID4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.310 1.505 0.690 ;
        RECT  1.450 1.110 1.505 1.490 ;
        RECT  1.150 0.310 1.450 1.490 ;
        RECT  0.840 0.310 1.150 0.690 ;
        RECT  0.840 1.110 1.150 1.490 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.240 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.690 ;
        RECT  0.185 -0.165 1.615 0.165 ;
        RECT  0.075 -0.165 0.185 0.590 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.110 1.725 1.965 ;
        RECT  0.725 1.635 1.615 1.965 ;
        RECT  0.535 1.410 0.725 1.965 ;
        RECT  0.000 1.635 0.535 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.840 0.310 1.050 0.690 ;
        RECT  0.840 1.110 1.050 1.490 ;
        RECT  0.730 0.780 0.940 0.890 ;
        RECT  0.640 0.480 0.730 1.320 ;
        RECT  0.295 0.480 0.640 0.590 ;
        RECT  0.185 1.210 0.640 1.320 ;
        RECT  0.075 1.210 0.185 1.485 ;
    END
END ISOHID4

MACRO ISOHID8
    CLASS CORE ;
    FOREIGN ISOHID8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.325 3.505 0.700 ;
        RECT  2.850 1.100 3.505 1.475 ;
        RECT  2.350 0.325 2.850 1.475 ;
        RECT  1.850 0.325 2.350 0.700 ;
        RECT  1.850 1.100 2.350 1.475 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.700 1.550 1.130 ;
        RECT  0.750 1.030 1.440 1.130 ;
        RECT  0.650 0.780 0.750 1.130 ;
        RECT  0.560 0.780 0.650 0.890 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.1646 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.600 1.150 0.920 ;
        RECT  0.170 0.600 1.040 0.690 ;
        RECT  0.050 0.600 0.170 1.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.165 3.800 0.165 ;
        RECT  3.615 -0.165 3.725 0.690 ;
        RECT  0.185 -0.165 3.615 0.165 ;
        RECT  0.075 -0.165 0.185 0.475 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 1.635 3.800 1.965 ;
        RECT  3.615 1.100 3.725 1.965 ;
        RECT  0.000 1.635 3.615 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.325 3.505 0.700 ;
        RECT  2.950 1.100 3.505 1.475 ;
        RECT  1.850 0.325 2.250 0.700 ;
        RECT  1.850 1.100 2.250 1.475 ;
        RECT  3.140 0.800 3.570 0.910 ;
        RECT  1.740 0.800 2.170 0.910 ;
        RECT  1.650 0.400 1.740 1.350 ;
        RECT  0.295 0.400 1.650 0.510 ;
        RECT  0.185 1.240 1.650 1.350 ;
        RECT  0.075 1.240 0.185 1.470 ;
    END
END ISOHID8

MACRO ISOLOD1
    CLASS CORE ;
    FOREIGN ISOLOD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.220 0.310 1.350 1.490 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.710 0.760 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.045 1.635 1.400 1.965 ;
        RECT  0.855 1.400 1.045 1.965 ;
        RECT  0.000 1.635 0.855 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.490 1.110 1.290 ;
        RECT  0.725 0.490 1.000 0.600 ;
        RECT  0.685 1.200 1.000 1.290 ;
        RECT  0.575 1.200 0.685 1.440 ;
        RECT  0.465 0.750 0.535 0.920 ;
        RECT  0.375 0.490 0.465 1.310 ;
        RECT  0.045 0.490 0.375 0.600 ;
        RECT  0.045 1.200 0.375 1.310 ;
    END
END ISOLOD1

MACRO ISOLOD2
    CLASS CORE ;
    FOREIGN ISOLOD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.455 0.555 1.550 1.245 ;
        RECT  1.450 0.310 1.455 1.490 ;
        RECT  1.345 0.310 1.450 0.690 ;
        RECT  1.345 1.110 1.450 1.490 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.780 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 -0.165 1.800 0.165 ;
        RECT  1.605 -0.165 1.715 0.445 ;
        RECT  1.235 -0.165 1.605 0.165 ;
        RECT  1.045 -0.165 1.235 0.410 ;
        RECT  0.000 -0.165 1.045 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.635 1.800 1.965 ;
        RECT  1.605 1.355 1.715 1.965 ;
        RECT  1.150 1.635 1.605 1.965 ;
        RECT  1.150 1.400 1.235 1.500 ;
        RECT  1.050 1.400 1.150 1.965 ;
        RECT  0.815 1.400 1.050 1.500 ;
        RECT  0.000 1.635 1.050 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.125 0.510 1.235 1.290 ;
        RECT  0.795 0.510 1.125 0.600 ;
        RECT  0.705 1.200 1.125 1.290 ;
        RECT  0.595 1.200 0.705 1.440 ;
        RECT  0.465 0.750 0.535 0.920 ;
        RECT  0.375 0.490 0.465 1.310 ;
        RECT  0.045 0.490 0.375 0.600 ;
        RECT  0.045 1.200 0.375 1.310 ;
    END
END ISOLOD2

MACRO ISOLOD4
    CLASS CORE ;
    FOREIGN ISOLOD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.310 1.905 0.690 ;
        RECT  1.850 1.110 1.905 1.490 ;
        RECT  1.550 0.310 1.850 1.490 ;
        RECT  1.240 0.310 1.550 0.690 ;
        RECT  1.240 1.110 1.550 1.490 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.710 0.760 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 -0.165 2.200 0.165 ;
        RECT  2.015 -0.165 2.125 0.690 ;
        RECT  0.000 -0.165 2.015 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 1.635 2.200 1.965 ;
        RECT  2.015 1.110 2.125 1.965 ;
        RECT  1.055 1.635 2.015 1.965 ;
        RECT  0.865 1.400 1.055 1.965 ;
        RECT  0.000 1.635 0.865 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.310 1.450 0.690 ;
        RECT  1.240 1.110 1.450 1.490 ;
        RECT  1.020 0.490 1.130 1.290 ;
        RECT  0.745 0.490 1.020 0.600 ;
        RECT  0.685 1.200 1.020 1.290 ;
        RECT  0.575 1.200 0.685 1.440 ;
        RECT  0.465 0.750 0.535 0.920 ;
        RECT  0.375 0.490 0.465 1.310 ;
        RECT  0.045 0.490 0.375 0.600 ;
        RECT  0.045 1.200 0.375 1.310 ;
    END
END ISOLOD4

MACRO ISOLOD8
    CLASS CORE ;
    FOREIGN ISOLOD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.325 3.905 0.700 ;
        RECT  3.250 1.100 3.905 1.475 ;
        RECT  2.750 0.325 3.250 1.475 ;
        RECT  2.250 0.325 2.750 0.700 ;
        RECT  2.250 1.100 2.750 1.475 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.700 1.950 1.120 ;
        RECT  0.955 1.020 1.840 1.120 ;
        RECT  0.845 0.750 0.955 1.120 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.690 ;
        RECT  0.485 -0.165 4.015 0.165 ;
        RECT  0.295 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.110 4.125 1.965 ;
        RECT  2.085 1.635 4.015 1.965 ;
        RECT  1.895 1.395 2.085 1.965 ;
        RECT  0.750 1.635 1.895 1.965 ;
        RECT  0.750 1.395 1.005 1.495 ;
        RECT  0.650 1.395 0.750 1.965 ;
        RECT  0.295 1.395 0.650 1.495 ;
        RECT  0.000 1.635 0.650 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.350 0.325 3.905 0.700 ;
        RECT  3.350 1.100 3.905 1.475 ;
        RECT  2.250 0.325 2.650 0.700 ;
        RECT  2.250 1.100 2.650 1.475 ;
        RECT  3.530 0.800 3.970 0.910 ;
        RECT  2.140 0.800 2.590 0.910 ;
        RECT  2.050 0.345 2.140 1.305 ;
        RECT  0.785 0.345 2.050 0.455 ;
        RECT  0.555 1.215 2.050 1.305 ;
        RECT  1.410 0.780 1.500 0.890 ;
        RECT  1.300 0.570 1.410 0.890 ;
        RECT  0.735 0.570 1.300 0.660 ;
        RECT  0.645 0.570 0.735 0.905 ;
        RECT  0.445 0.795 0.645 0.905 ;
        RECT  0.355 0.510 0.445 1.305 ;
        RECT  0.185 0.510 0.355 0.600 ;
        RECT  0.185 1.215 0.355 1.305 ;
        RECT  0.075 0.360 0.185 0.600 ;
        RECT  0.075 1.215 0.185 1.455 ;
    END
END ISOLOD8

MACRO LHCND1
    CLASS CORE ;
    FOREIGN LHCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1350 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.025 3.065 1.125 ;
        RECT  2.950 0.480 3.055 0.650 ;
        RECT  2.850 0.480 2.950 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.425 0.285 3.550 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.980 1.710 1.085 ;
        RECT  1.150 0.675 1.245 0.785 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.355 1.000 1.050 1.090 ;
        RECT  0.245 0.710 0.355 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.635 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.675 0.495 1.450 0.585 ;
        RECT  0.575 0.275 0.675 0.585 ;
        RECT  0.480 0.275 0.575 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 -0.165 3.600 0.165 ;
        RECT  3.100 -0.165 3.270 0.360 ;
        RECT  2.760 -0.165 3.100 0.165 ;
        RECT  2.660 -0.165 2.760 0.685 ;
        RECT  0.390 -0.165 2.660 0.165 ;
        RECT  0.390 0.495 0.485 0.585 ;
        RECT  0.290 -0.165 0.390 0.585 ;
        RECT  0.000 -0.165 0.290 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.635 3.600 1.965 ;
        RECT  3.100 1.415 3.270 1.965 ;
        RECT  2.805 1.635 3.100 1.965 ;
        RECT  2.615 1.395 2.805 1.965 ;
        RECT  0.000 1.635 2.615 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.175 0.740 3.295 1.305 ;
        RECT  2.570 1.215 3.175 1.305 ;
        RECT  2.500 0.305 2.570 1.305 ;
        RECT  2.470 0.305 2.500 1.465 ;
        RECT  2.355 0.305 2.470 0.405 ;
        RECT  2.400 1.215 2.470 1.465 ;
        RECT  2.280 0.740 2.380 0.930 ;
        RECT  2.190 0.515 2.280 1.495 ;
        RECT  1.680 1.395 2.190 1.495 ;
        RECT  2.000 0.315 2.100 1.275 ;
        RECT  1.125 0.315 2.000 0.405 ;
        RECT  1.285 1.175 2.000 1.275 ;
        RECT  0.185 1.405 1.420 1.505 ;
        RECT  0.540 1.180 1.285 1.275 ;
        RECT  0.155 1.255 0.185 1.505 ;
        RECT  0.155 0.405 0.180 0.600 ;
        RECT  0.065 0.405 0.155 1.505 ;
    END
END LHCND1

MACRO LHCND2
    CLASS CORE ;
    FOREIGN LHCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.275 2.960 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.465 0.510 3.550 1.195 ;
        RECT  3.450 0.275 3.465 1.490 ;
        RECT  3.355 0.275 3.450 0.675 ;
        RECT  3.355 1.045 3.450 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0810 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.000 1.750 1.105 ;
        RECT  1.150 0.675 1.240 0.785 ;
        RECT  1.050 0.675 1.150 1.105 ;
        RECT  0.355 1.000 1.050 1.105 ;
        RECT  0.240 0.700 0.355 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0406 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.495 1.875 0.660 ;
        RECT  1.445 0.495 1.555 0.890 ;
        RECT  0.650 0.495 1.445 0.585 ;
        RECT  0.550 0.275 0.650 0.585 ;
        RECT  0.445 0.275 0.550 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 -0.165 3.800 0.165 ;
        RECT  3.620 -0.165 3.720 0.445 ;
        RECT  0.000 -0.165 3.620 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.635 3.800 1.965 ;
        RECT  3.610 1.325 3.730 1.965 ;
        RECT  0.000 1.635 3.610 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.210 0.785 3.360 0.885 ;
        RECT  3.110 0.785 3.210 1.505 ;
        RECT  2.555 1.395 3.110 1.505 ;
        RECT  2.455 0.305 2.555 1.505 ;
        RECT  2.300 0.305 2.455 0.415 ;
        RECT  2.365 1.315 2.455 1.505 ;
        RECT  2.255 0.505 2.340 1.215 ;
        RECT  2.240 0.505 2.255 1.525 ;
        RECT  2.145 0.505 2.240 0.685 ;
        RECT  2.145 1.035 2.240 1.525 ;
        RECT  1.660 1.415 2.145 1.525 ;
        RECT  2.055 0.775 2.100 0.945 ;
        RECT  1.965 0.315 2.055 1.285 ;
        RECT  1.105 0.315 1.965 0.405 ;
        RECT  0.505 1.195 1.965 1.285 ;
        RECT  0.185 1.415 1.400 1.525 ;
        RECT  0.150 1.215 0.185 1.525 ;
        RECT  0.150 0.390 0.180 0.585 ;
        RECT  0.060 0.390 0.150 1.525 ;
    END
END LHCND2

MACRO LHCND4
    CLASS CORE ;
    FOREIGN LHCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.310 3.845 0.690 ;
        RECT  3.650 1.110 3.845 1.290 ;
        RECT  3.350 0.310 3.650 1.290 ;
        RECT  3.135 0.310 3.350 0.690 ;
        RECT  3.135 1.110 3.350 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.310 4.885 0.690 ;
        RECT  4.850 1.110 4.885 1.490 ;
        RECT  4.550 0.310 4.850 1.490 ;
        RECT  4.175 0.310 4.550 0.690 ;
        RECT  4.175 1.110 4.550 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0810 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.000 1.750 1.105 ;
        RECT  1.150 0.675 1.240 0.785 ;
        RECT  1.050 0.675 1.150 1.105 ;
        RECT  0.355 1.000 1.050 1.105 ;
        RECT  0.240 0.700 0.355 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0406 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.495 1.875 0.665 ;
        RECT  1.445 0.495 1.555 0.890 ;
        RECT  0.650 0.495 1.445 0.585 ;
        RECT  0.550 0.275 0.650 0.585 ;
        RECT  0.445 0.275 0.550 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 -0.165 5.200 0.165 ;
        RECT  4.995 -0.165 5.105 0.690 ;
        RECT  4.065 -0.165 4.995 0.165 ;
        RECT  3.955 -0.165 4.065 0.690 ;
        RECT  3.025 -0.165 3.955 0.165 ;
        RECT  2.915 -0.165 3.025 0.465 ;
        RECT  2.505 -0.165 2.915 0.165 ;
        RECT  2.395 -0.165 2.505 0.465 ;
        RECT  0.000 -0.165 2.395 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 1.635 5.200 1.965 ;
        RECT  4.995 1.110 5.105 1.965 ;
        RECT  2.505 1.635 4.995 1.965 ;
        RECT  2.395 1.305 2.505 1.965 ;
        RECT  0.000 1.635 2.395 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.175 0.310 4.450 0.690 ;
        RECT  4.175 1.110 4.450 1.490 ;
        RECT  3.750 0.310 3.845 0.690 ;
        RECT  3.750 1.110 3.845 1.290 ;
        RECT  3.135 0.310 3.250 0.690 ;
        RECT  3.135 1.110 3.250 1.290 ;
        RECT  4.065 0.800 4.320 0.900 ;
        RECT  3.955 0.800 4.065 1.525 ;
        RECT  2.875 1.415 3.955 1.525 ;
        RECT  2.765 0.555 2.875 1.525 ;
        RECT  2.655 0.310 2.765 0.690 ;
        RECT  2.655 1.110 2.765 1.525 ;
        RECT  2.340 0.800 2.660 0.900 ;
        RECT  2.255 0.555 2.340 1.210 ;
        RECT  2.240 0.310 2.255 1.525 ;
        RECT  2.145 0.310 2.240 0.685 ;
        RECT  2.145 1.110 2.240 1.525 ;
        RECT  1.670 1.415 2.145 1.525 ;
        RECT  2.055 0.775 2.100 0.945 ;
        RECT  1.965 0.315 2.055 1.285 ;
        RECT  1.125 0.315 1.965 0.405 ;
        RECT  0.515 1.195 1.965 1.285 ;
        RECT  0.185 1.415 1.390 1.525 ;
        RECT  0.150 1.215 0.185 1.525 ;
        RECT  0.150 0.390 0.180 0.585 ;
        RECT  0.060 0.390 0.150 1.525 ;
    END
END LHCND4

MACRO LHCNDD1
    CLASS CORE ;
    FOREIGN LHCNDD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1210 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.525 3.310 0.635 ;
        RECT  3.150 1.020 3.310 1.130 ;
        RECT  3.050 0.525 3.150 1.130 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.275 3.750 1.490 ;
        RECT  3.615 0.275 3.650 0.685 ;
        RECT  3.615 1.080 3.650 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.800 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.415 0.305 3.525 1.340 ;
        RECT  2.610 0.305 3.415 0.415 ;
        RECT  2.770 1.240 3.415 1.340 ;
        RECT  2.585 0.780 2.940 0.890 ;
        RECT  2.660 1.240 2.770 1.525 ;
        RECT  2.565 0.505 2.585 0.890 ;
        RECT  2.475 0.505 2.565 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.280 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.280 0.405 ;
        RECT  0.795 1.205 2.280 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCNDD1

MACRO LHCNDD2
    CLASS CORE ;
    FOREIGN LHCNDD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.525 3.350 1.130 ;
        RECT  3.150 0.525 3.250 0.635 ;
        RECT  3.150 1.020 3.250 1.130 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.585 3.950 1.180 ;
        RECT  3.830 0.585 3.850 0.685 ;
        RECT  3.830 1.080 3.850 1.180 ;
        RECT  3.720 0.275 3.830 0.685 ;
        RECT  3.720 1.080 3.830 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0419 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.090 -0.165 4.200 0.165 ;
        RECT  3.980 -0.165 4.090 0.485 ;
        RECT  0.000 -0.165 3.980 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.090 1.635 4.200 1.965 ;
        RECT  3.980 1.280 4.090 1.965 ;
        RECT  3.600 1.635 3.980 1.965 ;
        RECT  3.430 1.400 3.600 1.965 ;
        RECT  3.080 1.635 3.430 1.965 ;
        RECT  2.910 1.400 3.080 1.965 ;
        RECT  0.000 1.635 2.910 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.630 0.780 3.755 0.890 ;
        RECT  3.520 0.305 3.630 1.310 ;
        RECT  2.640 0.305 3.520 0.415 ;
        RECT  2.800 1.220 3.520 1.310 ;
        RECT  2.615 0.780 3.060 0.890 ;
        RECT  2.690 1.220 2.800 1.525 ;
        RECT  2.595 0.505 2.615 0.890 ;
        RECT  2.505 0.505 2.595 1.525 ;
        RECT  2.010 1.415 2.505 1.525 ;
        RECT  2.320 0.295 2.410 1.315 ;
        RECT  1.465 0.295 2.320 0.405 ;
        RECT  0.795 1.205 2.320 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCNDD2

MACRO LHCNDD4
    CLASS CORE ;
    FOREIGN LHCNDD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.325 4.125 0.635 ;
        RECT  3.850 1.110 4.085 1.290 ;
        RECT  3.550 0.325 3.850 1.290 ;
        RECT  3.415 0.325 3.550 0.635 ;
        RECT  3.455 1.110 3.550 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.325 5.150 0.635 ;
        RECT  5.050 1.100 5.150 1.410 ;
        RECT  4.750 0.325 5.050 1.410 ;
        RECT  4.415 0.325 4.750 0.635 ;
        RECT  4.415 1.100 4.750 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.415 0.325 4.650 0.635 ;
        RECT  4.415 1.100 4.650 1.410 ;
        RECT  3.950 0.325 4.125 0.635 ;
        RECT  3.950 1.110 4.085 1.290 ;
        RECT  3.415 0.325 3.450 0.635 ;
        RECT  4.295 0.780 4.500 0.890 ;
        RECT  4.195 0.780 4.295 1.480 ;
        RECT  3.290 1.380 4.195 1.480 ;
        RECT  3.200 0.575 3.290 1.480 ;
        RECT  3.075 0.575 3.200 0.685 ;
        RECT  3.075 1.380 3.200 1.480 ;
        RECT  2.965 0.275 3.075 0.685 ;
        RECT  2.965 1.050 3.075 1.480 ;
        RECT  2.585 0.780 3.050 0.890 ;
        RECT  2.475 0.275 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.290 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.290 0.405 ;
        RECT  0.795 1.205 2.290 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCNDD4

MACRO LHCNDQD1
    CLASS CORE ;
    FOREIGN LHCNDQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.275 3.350 1.490 ;
        RECT  3.215 0.275 3.250 0.675 ;
        RECT  3.215 1.080 3.250 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0469 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.100 0.495 2.210 0.690 ;
        RECT  0.950 0.495 2.100 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.065 -0.165 3.400 0.165 ;
        RECT  2.955 -0.165 3.065 0.485 ;
        RECT  0.880 -0.165 2.955 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.065 1.635 3.400 1.965 ;
        RECT  2.955 1.280 3.065 1.965 ;
        RECT  0.000 1.635 2.955 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.120 0.750 3.160 0.920 ;
        RECT  3.030 0.575 3.120 1.180 ;
        RECT  2.805 0.575 3.030 0.675 ;
        RECT  2.805 1.080 3.030 1.180 ;
        RECT  2.605 0.780 2.940 0.890 ;
        RECT  2.695 0.255 2.805 0.675 ;
        RECT  2.695 1.080 2.805 1.525 ;
        RECT  2.505 0.505 2.605 1.525 ;
        RECT  2.040 1.415 2.505 1.525 ;
        RECT  2.310 0.295 2.410 1.315 ;
        RECT  1.505 0.295 2.310 0.405 ;
        RECT  0.795 1.205 2.310 1.315 ;
        RECT  1.580 0.995 2.060 1.105 ;
        RECT  1.575 1.435 1.785 1.545 ;
        RECT  1.470 0.675 1.580 1.105 ;
        RECT  0.460 1.435 1.575 1.525 ;
        RECT  0.700 1.010 1.470 1.105 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCNDQD1

MACRO LHCNDQD2
    CLASS CORE ;
    FOREIGN LHCNDQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.590 3.550 1.180 ;
        RECT  3.350 0.590 3.450 0.690 ;
        RECT  3.350 1.080 3.450 1.180 ;
        RECT  3.165 0.275 3.350 0.690 ;
        RECT  3.165 1.080 3.350 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.075 0.780 3.300 0.890 ;
        RECT  2.975 0.305 3.075 1.310 ;
        RECT  2.625 0.305 2.975 0.415 ;
        RECT  2.775 1.220 2.975 1.310 ;
        RECT  2.585 0.780 2.875 0.890 ;
        RECT  2.665 1.220 2.775 1.525 ;
        RECT  2.575 0.505 2.585 0.890 ;
        RECT  2.475 0.505 2.575 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.290 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.290 0.405 ;
        RECT  0.795 1.205 2.290 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCNDQD2

MACRO LHCNDQD4
    CLASS CORE ;
    FOREIGN LHCNDQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.325 4.150 0.635 ;
        RECT  4.050 1.100 4.150 1.410 ;
        RECT  3.750 0.325 4.050 1.410 ;
        RECT  3.415 0.325 3.750 0.635 ;
        RECT  3.415 1.100 3.750 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.415 0.325 3.650 0.635 ;
        RECT  3.415 1.100 3.650 1.410 ;
        RECT  3.290 0.780 3.600 0.890 ;
        RECT  3.190 0.575 3.290 1.150 ;
        RECT  3.075 0.575 3.190 0.685 ;
        RECT  3.075 1.050 3.190 1.150 ;
        RECT  2.595 0.780 3.080 0.890 ;
        RECT  2.965 0.275 3.075 0.685 ;
        RECT  2.965 1.050 3.075 1.460 ;
        RECT  2.495 0.275 2.595 1.525 ;
        RECT  2.010 1.415 2.495 1.525 ;
        RECT  2.310 0.295 2.400 1.315 ;
        RECT  1.465 0.295 2.310 0.405 ;
        RECT  0.795 1.205 2.310 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCNDQD4

MACRO LHCNQD1
    CLASS CORE ;
    FOREIGN LHCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.150 1.490 ;
        RECT  3.015 0.275 3.050 0.665 ;
        RECT  3.015 1.040 3.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.185 1.015 1.775 1.105 ;
        RECT  1.185 0.645 1.280 0.755 ;
        RECT  1.075 0.645 1.185 1.105 ;
        RECT  0.350 1.015 1.075 1.105 ;
        RECT  0.250 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0421 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.965 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0413 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 0.465 1.950 0.735 ;
        RECT  1.550 0.465 1.820 0.555 ;
        RECT  1.435 0.465 1.550 0.890 ;
        RECT  0.750 0.465 1.435 0.555 ;
        RECT  0.650 0.255 0.750 0.555 ;
        RECT  0.475 0.255 0.650 0.345 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.865 -0.165 3.200 0.165 ;
        RECT  2.755 -0.165 2.865 0.660 ;
        RECT  0.365 -0.165 2.755 0.165 ;
        RECT  0.365 0.480 0.495 0.590 ;
        RECT  0.275 -0.165 0.365 0.590 ;
        RECT  0.000 -0.165 0.275 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.865 1.635 3.200 1.965 ;
        RECT  2.755 1.040 2.865 1.965 ;
        RECT  0.000 1.635 2.755 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.635 0.750 2.950 0.920 ;
        RECT  2.535 0.255 2.635 1.225 ;
        RECT  2.420 0.255 2.535 0.365 ;
        RECT  2.495 1.015 2.535 1.225 ;
        RECT  2.385 0.735 2.435 0.945 ;
        RECT  2.365 0.735 2.385 1.505 ;
        RECT  2.265 0.480 2.365 1.505 ;
        RECT  1.750 1.395 2.265 1.505 ;
        RECT  2.075 0.275 2.175 1.285 ;
        RECT  1.170 0.275 2.075 0.375 ;
        RECT  0.525 1.195 2.075 1.285 ;
        RECT  1.260 1.395 1.470 1.505 ;
        RECT  0.185 1.395 1.260 1.485 ;
        RECT  0.160 0.385 0.185 0.590 ;
        RECT  0.160 1.255 0.185 1.485 ;
        RECT  0.060 0.385 0.160 1.485 ;
    END
END LHCNQD1

MACRO LHCNQD2
    CLASS CORE ;
    FOREIGN LHCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.150 1.490 ;
        RECT  2.965 0.275 3.050 0.665 ;
        RECT  2.965 1.040 3.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.185 1.015 1.770 1.105 ;
        RECT  1.185 0.645 1.280 0.755 ;
        RECT  1.075 0.645 1.185 1.105 ;
        RECT  0.350 1.015 1.075 1.105 ;
        RECT  0.250 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0421 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.965 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0415 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 0.465 1.950 0.735 ;
        RECT  1.550 0.465 1.820 0.555 ;
        RECT  1.435 0.465 1.550 0.890 ;
        RECT  0.750 0.465 1.435 0.555 ;
        RECT  0.650 0.255 0.750 0.555 ;
        RECT  0.475 0.255 0.650 0.345 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.365 -0.165 3.400 0.165 ;
        RECT  0.365 0.480 0.495 0.590 ;
        RECT  0.275 -0.165 0.365 0.590 ;
        RECT  0.000 -0.165 0.275 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.635 0.780 2.950 0.890 ;
        RECT  2.535 0.305 2.635 1.175 ;
        RECT  2.415 0.305 2.535 0.415 ;
        RECT  2.430 1.065 2.535 1.175 ;
        RECT  2.350 0.735 2.435 0.945 ;
        RECT  2.340 1.395 2.385 1.505 ;
        RECT  2.340 0.495 2.350 0.945 ;
        RECT  2.250 0.495 2.340 1.505 ;
        RECT  1.740 1.395 2.250 1.505 ;
        RECT  2.060 0.275 2.160 1.285 ;
        RECT  1.170 0.275 2.060 0.375 ;
        RECT  0.525 1.195 2.060 1.285 ;
        RECT  1.260 1.395 1.470 1.505 ;
        RECT  0.185 1.395 1.260 1.485 ;
        RECT  0.160 0.355 0.185 0.565 ;
        RECT  0.160 1.215 0.185 1.485 ;
        RECT  0.060 0.355 0.160 1.485 ;
    END
END LHCNQD2

MACRO LHCNQD4
    CLASS CORE ;
    FOREIGN LHCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 0.310 3.860 0.690 ;
        RECT  3.750 1.110 3.860 1.490 ;
        RECT  3.650 0.545 3.750 0.690 ;
        RECT  3.650 1.110 3.750 1.210 ;
        RECT  3.350 0.545 3.650 1.210 ;
        RECT  3.240 0.310 3.350 0.690 ;
        RECT  3.345 1.110 3.350 1.210 ;
        RECT  3.240 1.110 3.345 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.185 1.015 1.770 1.105 ;
        RECT  1.185 0.645 1.280 0.755 ;
        RECT  1.075 0.645 1.185 1.105 ;
        RECT  0.350 1.015 1.075 1.105 ;
        RECT  0.250 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0421 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.965 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0415 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 0.465 1.950 0.735 ;
        RECT  1.550 0.465 1.820 0.555 ;
        RECT  1.435 0.465 1.550 0.890 ;
        RECT  0.750 0.465 1.435 0.555 ;
        RECT  0.650 0.255 0.750 0.555 ;
        RECT  0.475 0.255 0.650 0.345 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.690 ;
        RECT  3.605 -0.165 4.015 0.165 ;
        RECT  3.495 -0.165 3.605 0.455 ;
        RECT  3.085 -0.165 3.495 0.165 ;
        RECT  2.975 -0.165 3.085 0.690 ;
        RECT  0.365 -0.165 2.975 0.165 ;
        RECT  0.365 0.480 0.495 0.590 ;
        RECT  0.275 -0.165 0.365 0.590 ;
        RECT  0.000 -0.165 0.275 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.110 4.125 1.965 ;
        RECT  3.605 1.635 4.015 1.965 ;
        RECT  3.495 1.320 3.605 1.965 ;
        RECT  3.085 1.635 3.495 1.965 ;
        RECT  2.975 1.110 3.085 1.965 ;
        RECT  0.000 1.635 2.975 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 0.310 3.860 0.690 ;
        RECT  3.750 1.110 3.860 1.490 ;
        RECT  3.240 0.310 3.250 0.690 ;
        RECT  3.240 1.110 3.250 1.490 ;
        RECT  2.825 0.800 3.260 0.910 ;
        RECT  2.715 0.310 2.825 1.490 ;
        RECT  2.350 0.800 2.560 0.910 ;
        RECT  2.350 1.395 2.385 1.505 ;
        RECT  2.250 0.495 2.350 1.505 ;
        RECT  1.740 1.395 2.250 1.505 ;
        RECT  2.060 0.275 2.160 1.285 ;
        RECT  1.170 0.275 2.060 0.375 ;
        RECT  0.525 1.195 2.060 1.285 ;
        RECT  1.260 1.395 1.470 1.505 ;
        RECT  0.185 1.395 1.260 1.485 ;
        RECT  0.160 0.355 0.185 0.565 ;
        RECT  0.160 1.215 0.185 1.485 ;
        RECT  0.060 0.355 0.160 1.485 ;
    END
END LHCNQD4

MACRO LHCSND1
    CLASS CORE ;
    FOREIGN LHCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.370 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.500 3.245 0.675 ;
        RECT  3.150 1.025 3.245 1.125 ;
        RECT  3.050 0.500 3.150 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.275 3.750 1.490 ;
        RECT  3.625 0.275 3.650 0.695 ;
        RECT  3.615 1.040 3.650 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.980 1.725 1.090 ;
        RECT  1.150 0.675 1.270 0.775 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.350 1.000 1.050 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0411 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.435 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.435 0.585 ;
        RECT  0.650 0.255 0.750 0.585 ;
        RECT  0.480 0.255 0.650 0.365 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 -0.165 3.800 0.165 ;
        RECT  3.355 -0.165 3.465 0.585 ;
        RECT  2.690 -0.165 3.355 0.165 ;
        RECT  2.550 -0.165 2.690 0.375 ;
        RECT  0.385 -0.165 2.550 0.165 ;
        RECT  0.385 0.475 0.495 0.585 ;
        RECT  0.285 -0.165 0.385 0.585 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.495 1.635 3.800 1.965 ;
        RECT  3.325 1.395 3.495 1.965 ;
        RECT  2.655 1.635 3.325 1.965 ;
        RECT  2.445 1.390 2.655 1.965 ;
        RECT  0.000 1.635 2.445 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.460 0.730 3.540 0.940 ;
        RECT  3.360 0.730 3.460 1.305 ;
        RECT  2.930 1.215 3.360 1.305 ;
        RECT  2.930 0.305 3.025 0.410 ;
        RECT  2.820 0.305 2.930 1.470 ;
        RECT  2.610 0.490 2.720 1.300 ;
        RECT  2.315 0.490 2.610 0.600 ;
        RECT  2.295 1.200 2.610 1.300 ;
        RECT  2.185 1.200 2.295 1.505 ;
        RECT  1.695 1.395 2.185 1.505 ;
        RECT  2.095 0.315 2.120 0.930 ;
        RECT  2.000 0.315 2.095 1.285 ;
        RECT  1.145 0.315 2.000 0.405 ;
        RECT  0.520 1.180 2.000 1.285 ;
        RECT  0.185 1.395 1.405 1.505 ;
        RECT  0.160 0.385 0.185 0.585 ;
        RECT  0.160 1.255 0.185 1.505 ;
        RECT  0.060 0.385 0.160 1.505 ;
    END
END LHCSND1

MACRO LHCSND2
    CLASS CORE ;
    FOREIGN LHCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.710 2.550 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 1.025 3.395 1.125 ;
        RECT  3.230 0.275 3.350 1.125 ;
        RECT  3.185 1.025 3.230 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.865 0.510 3.950 1.100 ;
        RECT  3.850 0.275 3.865 1.490 ;
        RECT  3.755 0.275 3.850 0.695 ;
        RECT  3.755 0.995 3.850 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0802 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.980 1.725 1.090 ;
        RECT  1.150 0.675 1.270 0.775 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.350 1.000 1.050 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0415 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.435 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.435 0.585 ;
        RECT  0.650 0.255 0.750 0.585 ;
        RECT  0.480 0.255 0.650 0.365 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.445 ;
        RECT  3.605 -0.165 4.015 0.165 ;
        RECT  3.495 -0.165 3.605 0.695 ;
        RECT  0.385 -0.165 3.495 0.165 ;
        RECT  0.385 0.475 0.495 0.585 ;
        RECT  0.285 -0.165 0.385 0.585 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.210 4.125 1.965 ;
        RECT  3.360 1.635 4.015 1.965 ;
        RECT  3.360 1.395 3.645 1.505 ;
        RECT  3.220 1.395 3.360 1.965 ;
        RECT  2.935 1.395 3.220 1.505 ;
        RECT  2.555 1.635 3.220 1.965 ;
        RECT  2.445 1.200 2.555 1.965 ;
        RECT  0.000 1.635 2.445 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.615 0.785 3.740 0.890 ;
        RECT  3.505 0.785 3.615 1.305 ;
        RECT  2.825 1.215 3.505 1.305 ;
        RECT  2.935 0.330 3.065 0.940 ;
        RECT  2.345 0.330 2.935 0.445 ;
        RECT  2.715 0.545 2.825 1.470 ;
        RECT  2.625 0.545 2.715 0.650 ;
        RECT  2.235 0.330 2.345 1.505 ;
        RECT  1.695 1.395 2.235 1.505 ;
        RECT  2.015 0.315 2.125 1.285 ;
        RECT  1.145 0.315 2.015 0.405 ;
        RECT  0.520 1.180 2.015 1.285 ;
        RECT  0.185 1.395 1.405 1.505 ;
        RECT  0.160 0.390 0.185 0.580 ;
        RECT  0.160 1.195 0.185 1.505 ;
        RECT  0.060 0.390 0.160 1.505 ;
    END
END LHCSND2

MACRO LHCSND4
    CLASS CORE ;
    FOREIGN LHCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.700 2.550 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.310 4.315 0.695 ;
        RECT  4.050 1.110 4.315 1.290 ;
        RECT  3.750 0.310 4.050 1.290 ;
        RECT  3.625 0.310 3.750 0.695 ;
        RECT  3.625 1.110 3.750 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.310 5.350 0.690 ;
        RECT  5.250 1.110 5.350 1.490 ;
        RECT  4.950 0.310 5.250 1.490 ;
        RECT  4.625 0.310 4.950 0.690 ;
        RECT  4.625 1.110 4.950 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0802 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.980 1.720 1.090 ;
        RECT  1.150 0.675 1.270 0.775 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.350 1.000 1.050 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0415 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.435 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.435 0.585 ;
        RECT  0.650 0.255 0.750 0.585 ;
        RECT  0.480 0.255 0.650 0.365 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.385 -0.165 5.600 0.165 ;
        RECT  0.385 0.475 0.495 0.585 ;
        RECT  0.285 -0.165 0.385 0.585 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.625 0.310 4.850 0.690 ;
        RECT  4.625 1.110 4.850 1.490 ;
        RECT  4.150 0.310 4.315 0.695 ;
        RECT  4.150 1.110 4.315 1.290 ;
        RECT  3.625 0.310 3.650 0.695 ;
        RECT  3.625 1.110 3.650 1.290 ;
        RECT  4.515 0.800 4.760 0.910 ;
        RECT  4.425 0.800 4.515 1.505 ;
        RECT  3.275 1.400 4.425 1.505 ;
        RECT  3.380 0.600 3.490 1.200 ;
        RECT  3.275 0.600 3.380 0.690 ;
        RECT  3.275 1.110 3.380 1.200 ;
        RECT  3.165 0.310 3.275 0.690 ;
        RECT  3.165 1.110 3.275 1.505 ;
        RECT  3.075 0.800 3.270 0.910 ;
        RECT  2.965 0.345 3.075 1.505 ;
        RECT  2.365 0.345 2.965 0.455 ;
        RECT  1.690 1.395 2.965 1.505 ;
        RECT  2.745 0.700 2.855 1.285 ;
        RECT  2.120 1.180 2.745 1.285 ;
        RECT  2.010 0.315 2.120 1.285 ;
        RECT  1.145 0.315 2.010 0.405 ;
        RECT  0.520 1.180 2.010 1.285 ;
        RECT  0.185 1.395 1.410 1.505 ;
        RECT  0.160 0.390 0.185 0.580 ;
        RECT  0.160 1.195 0.185 1.505 ;
        RECT  0.060 0.390 0.160 1.505 ;
    END
END LHCSND4

MACRO LHCSNDD1
    CLASS CORE ;
    FOREIGN LHCSNDD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.750 1.090 ;
        RECT  2.630 0.710 2.650 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 1.015 3.655 1.125 ;
        RECT  3.550 0.275 3.605 0.675 ;
        RECT  3.450 0.275 3.550 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.275 4.150 1.490 ;
        RECT  4.025 0.275 4.050 0.675 ;
        RECT  4.015 1.080 4.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.865 -0.165 4.200 0.165 ;
        RECT  3.755 -0.165 3.865 0.655 ;
        RECT  3.070 -0.165 3.755 0.165 ;
        RECT  2.960 -0.165 3.070 0.355 ;
        RECT  0.880 -0.165 2.960 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.895 1.635 4.200 1.965 ;
        RECT  3.725 1.395 3.895 1.965 ;
        RECT  3.030 1.635 3.725 1.965 ;
        RECT  2.860 1.495 3.030 1.965 ;
        RECT  0.000 1.635 2.860 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.870 0.750 3.950 0.920 ;
        RECT  3.770 0.750 3.870 1.305 ;
        RECT  3.355 1.215 3.770 1.305 ;
        RECT  3.245 0.275 3.355 1.460 ;
        RECT  3.025 0.490 3.135 1.300 ;
        RECT  2.675 0.490 3.025 0.600 ;
        RECT  2.645 1.200 3.025 1.300 ;
        RECT  2.535 1.200 2.645 1.525 ;
        RECT  2.010 1.415 2.535 1.525 ;
        RECT  2.380 0.750 2.480 0.920 ;
        RECT  2.280 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.280 0.405 ;
        RECT  0.795 1.205 2.280 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCSNDD1

MACRO LHCSNDD2
    CLASS CORE ;
    FOREIGN LHCSNDD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.750 2.670 0.920 ;
        RECT  2.550 0.600 2.615 0.920 ;
        RECT  2.525 0.310 2.550 0.920 ;
        RECT  2.450 0.310 2.525 0.690 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.275 3.565 1.180 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.065 0.585 4.150 1.150 ;
        RECT  4.050 0.275 4.065 1.460 ;
        RECT  3.955 0.275 4.050 0.685 ;
        RECT  3.955 1.050 4.050 1.460 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.485 ;
        RECT  0.000 -0.165 4.215 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.250 4.325 1.965 ;
        RECT  0.000 1.635 4.215 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.820 0.780 3.960 0.890 ;
        RECT  3.720 0.780 3.820 1.370 ;
        RECT  3.295 1.270 3.720 1.370 ;
        RECT  3.195 0.575 3.295 1.370 ;
        RECT  3.065 0.575 3.195 0.685 ;
        RECT  3.065 1.270 3.195 1.370 ;
        RECT  2.865 0.780 3.095 0.890 ;
        RECT  2.955 0.275 3.065 0.685 ;
        RECT  2.955 1.050 3.065 1.460 ;
        RECT  2.815 0.575 2.865 1.150 ;
        RECT  2.775 0.275 2.815 1.150 ;
        RECT  2.705 0.275 2.775 0.665 ;
        RECT  2.585 1.050 2.775 1.150 ;
        RECT  2.475 1.050 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.350 0.780 2.430 0.890 ;
        RECT  2.260 0.295 2.350 1.315 ;
        RECT  1.465 0.295 2.260 0.405 ;
        RECT  0.795 1.205 2.260 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCSNDD2

MACRO LHCSNDD4
    CLASS CORE ;
    FOREIGN LHCSNDD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.700 2.760 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.325 4.665 0.635 ;
        RECT  4.450 1.110 4.655 1.290 ;
        RECT  4.150 0.325 4.450 1.290 ;
        RECT  3.945 0.325 4.150 0.635 ;
        RECT  3.955 1.110 4.150 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.325 5.685 0.635 ;
        RECT  5.650 1.100 5.685 1.410 ;
        RECT  5.350 0.325 5.650 1.410 ;
        RECT  4.965 0.325 5.350 0.635 ;
        RECT  4.965 1.100 5.350 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.895 -0.165 6.000 0.165 ;
        RECT  5.785 -0.165 5.895 0.685 ;
        RECT  0.000 -0.165 5.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.895 1.635 6.000 1.965 ;
        RECT  5.785 1.050 5.895 1.965 ;
        RECT  0.000 1.635 5.785 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.965 0.325 5.250 0.635 ;
        RECT  4.965 1.100 5.250 1.410 ;
        RECT  4.550 0.325 4.665 0.635 ;
        RECT  4.550 1.110 4.655 1.290 ;
        RECT  3.945 0.325 4.050 0.635 ;
        RECT  3.955 1.110 4.050 1.290 ;
        RECT  4.865 0.780 5.110 0.890 ;
        RECT  4.775 0.780 4.865 1.505 ;
        RECT  3.595 1.400 4.775 1.505 ;
        RECT  3.735 0.600 3.835 1.195 ;
        RECT  3.595 0.600 3.735 0.690 ;
        RECT  3.595 1.095 3.735 1.195 ;
        RECT  3.485 0.310 3.595 0.690 ;
        RECT  3.485 1.095 3.595 1.505 ;
        RECT  3.395 0.780 3.590 0.890 ;
        RECT  3.295 0.490 3.395 1.495 ;
        RECT  2.675 0.490 3.295 0.600 ;
        RECT  2.525 1.385 3.295 1.495 ;
        RECT  3.070 0.750 3.180 1.285 ;
        RECT  2.420 1.180 3.070 1.285 ;
        RECT  2.415 1.385 2.525 1.525 ;
        RECT  2.310 0.295 2.420 1.285 ;
        RECT  2.010 1.415 2.415 1.525 ;
        RECT  1.465 0.295 2.310 0.405 ;
        RECT  2.230 1.180 2.310 1.285 ;
        RECT  2.130 1.180 2.230 1.315 ;
        RECT  0.795 1.205 2.130 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCSNDD4

MACRO LHCSNDQD1
    CLASS CORE ;
    FOREIGN LHCSNDQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.770 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.275 3.550 1.490 ;
        RECT  3.415 0.275 3.450 0.675 ;
        RECT  3.415 1.080 3.450 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.600 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.305 0.750 3.360 0.920 ;
        RECT  3.205 0.310 3.305 1.145 ;
        RECT  2.865 0.310 3.205 0.420 ;
        RECT  2.865 1.035 3.205 1.145 ;
        RECT  2.985 0.510 3.095 0.930 ;
        RECT  2.560 0.510 2.985 0.620 ;
        RECT  2.560 1.250 2.575 1.525 ;
        RECT  2.470 0.510 2.560 1.525 ;
        RECT  2.010 1.415 2.470 1.525 ;
        RECT  2.280 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.280 0.405 ;
        RECT  0.795 1.205 2.280 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCSNDQD1

MACRO LHCSNDQD2
    CLASS CORE ;
    FOREIGN LHCSNDQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.750 2.670 0.920 ;
        RECT  2.550 0.600 2.615 0.920 ;
        RECT  2.525 0.310 2.550 0.920 ;
        RECT  2.450 0.310 2.525 0.690 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.585 3.750 1.150 ;
        RECT  3.615 0.585 3.650 0.685 ;
        RECT  3.615 1.050 3.650 1.150 ;
        RECT  3.505 0.275 3.615 0.685 ;
        RECT  3.505 1.050 3.615 1.460 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.875 -0.165 4.000 0.165 ;
        RECT  3.765 -0.165 3.875 0.475 ;
        RECT  3.365 -0.165 3.765 0.165 ;
        RECT  3.245 -0.165 3.365 0.475 ;
        RECT  0.000 -0.165 3.245 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.875 1.635 4.000 1.965 ;
        RECT  3.765 1.250 3.875 1.965 ;
        RECT  3.365 1.635 3.765 1.965 ;
        RECT  3.245 1.250 3.365 1.965 ;
        RECT  2.845 1.635 3.245 1.965 ;
        RECT  2.735 1.250 2.845 1.965 ;
        RECT  0.000 1.635 2.735 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.325 0.780 3.540 0.890 ;
        RECT  3.225 0.575 3.325 1.150 ;
        RECT  3.095 0.575 3.225 0.685 ;
        RECT  3.095 1.050 3.225 1.150 ;
        RECT  2.865 0.780 3.125 0.890 ;
        RECT  2.985 0.275 3.095 0.685 ;
        RECT  2.985 1.050 3.095 1.460 ;
        RECT  2.815 0.575 2.865 1.150 ;
        RECT  2.775 0.275 2.815 1.150 ;
        RECT  2.705 0.275 2.775 0.665 ;
        RECT  2.585 1.050 2.775 1.150 ;
        RECT  2.475 1.050 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.350 0.780 2.430 0.890 ;
        RECT  2.260 0.295 2.350 1.315 ;
        RECT  1.465 0.295 2.260 0.405 ;
        RECT  0.795 1.205 2.260 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCSNDQD2

MACRO LHCSNDQD4
    CLASS CORE ;
    FOREIGN LHCSNDQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.750 1.090 ;
        RECT  2.570 0.710 2.650 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.325 4.350 0.635 ;
        RECT  4.250 1.100 4.350 1.410 ;
        RECT  3.950 0.325 4.250 1.410 ;
        RECT  3.615 0.325 3.950 0.635 ;
        RECT  3.615 1.100 3.950 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.960 1.635 4.600 1.965 ;
        RECT  2.790 1.390 2.960 1.965 ;
        RECT  0.000 1.635 2.790 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.615 0.325 3.850 0.635 ;
        RECT  3.615 1.100 3.850 1.410 ;
        RECT  3.505 0.780 3.770 0.890 ;
        RECT  3.405 0.575 3.505 1.150 ;
        RECT  3.275 0.575 3.405 0.685 ;
        RECT  3.275 1.050 3.405 1.150 ;
        RECT  2.960 0.780 3.305 0.890 ;
        RECT  3.165 0.275 3.275 0.685 ;
        RECT  3.165 1.050 3.275 1.460 ;
        RECT  2.860 0.490 2.960 1.300 ;
        RECT  2.635 0.490 2.860 0.600 ;
        RECT  2.585 1.200 2.860 1.300 ;
        RECT  2.475 1.200 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.350 0.750 2.420 0.920 ;
        RECT  2.260 0.295 2.350 1.315 ;
        RECT  1.465 0.295 2.260 0.405 ;
        RECT  0.795 1.205 2.260 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.460 1.435 1.535 1.525 ;
        RECT  0.700 1.010 1.440 1.105 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHCSNDQD4

MACRO LHCSNQD1
    CLASS CORE ;
    FOREIGN LHCSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.370 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.275 3.350 1.490 ;
        RECT  3.220 0.275 3.250 0.695 ;
        RECT  3.215 1.040 3.250 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.980 1.725 1.090 ;
        RECT  1.150 0.675 1.270 0.775 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.350 1.000 1.050 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0411 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.435 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.435 0.585 ;
        RECT  0.650 0.255 0.750 0.585 ;
        RECT  0.480 0.255 0.650 0.365 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.065 -0.165 3.400 0.165 ;
        RECT  2.955 -0.165 3.065 0.585 ;
        RECT  0.385 -0.165 2.955 0.165 ;
        RECT  0.385 0.475 0.495 0.585 ;
        RECT  0.285 -0.165 0.385 0.585 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.065 1.635 3.400 1.965 ;
        RECT  2.955 1.040 3.065 1.965 ;
        RECT  2.580 1.635 2.955 1.965 ;
        RECT  2.400 1.390 2.580 1.965 ;
        RECT  0.000 1.635 2.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.845 0.740 3.140 0.930 ;
        RECT  2.805 0.545 2.845 1.135 ;
        RECT  2.745 0.275 2.805 1.490 ;
        RECT  2.695 0.275 2.745 0.675 ;
        RECT  2.695 1.035 2.745 1.490 ;
        RECT  2.560 0.750 2.635 0.930 ;
        RECT  2.460 0.425 2.560 1.300 ;
        RECT  2.335 0.425 2.460 0.535 ;
        RECT  2.285 1.200 2.460 1.300 ;
        RECT  2.180 1.200 2.285 1.505 ;
        RECT  1.695 1.395 2.180 1.505 ;
        RECT  2.090 0.315 2.120 0.930 ;
        RECT  2.000 0.315 2.090 1.285 ;
        RECT  1.145 0.315 2.000 0.405 ;
        RECT  0.520 1.180 2.000 1.285 ;
        RECT  0.185 1.395 1.415 1.505 ;
        RECT  0.160 0.385 0.185 0.585 ;
        RECT  0.160 1.255 0.185 1.505 ;
        RECT  0.060 0.385 0.160 1.505 ;
    END
END LHCSNQD1

MACRO LHCSNQD2
    CLASS CORE ;
    FOREIGN LHCSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.370 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.265 0.510 3.350 1.100 ;
        RECT  3.260 0.510 3.265 1.490 ;
        RECT  3.250 0.285 3.260 1.490 ;
        RECT  3.160 0.285 3.250 0.675 ;
        RECT  3.155 1.000 3.250 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0802 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.980 1.725 1.090 ;
        RECT  1.150 0.675 1.270 0.775 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.350 1.000 1.050 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0415 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.435 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.435 0.585 ;
        RECT  0.650 0.255 0.750 0.585 ;
        RECT  0.480 0.255 0.650 0.365 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 -0.165 3.600 0.165 ;
        RECT  3.420 -0.165 3.525 0.445 ;
        RECT  3.005 -0.165 3.420 0.165 ;
        RECT  2.895 -0.165 3.005 0.495 ;
        RECT  0.385 -0.165 2.895 0.165 ;
        RECT  0.385 0.475 0.495 0.585 ;
        RECT  0.285 -0.165 0.385 0.585 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 1.635 3.600 1.965 ;
        RECT  3.415 1.210 3.525 1.965 ;
        RECT  2.595 1.635 3.415 1.965 ;
        RECT  2.395 1.390 2.595 1.965 ;
        RECT  0.000 1.635 2.395 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.000 0.785 3.140 0.890 ;
        RECT  2.900 0.585 3.000 1.095 ;
        RECT  2.745 0.585 2.900 0.695 ;
        RECT  2.765 0.995 2.900 1.095 ;
        RECT  2.550 0.785 2.790 0.890 ;
        RECT  2.655 0.995 2.765 1.245 ;
        RECT  2.640 0.275 2.745 0.695 ;
        RECT  2.460 0.425 2.550 1.300 ;
        RECT  2.325 0.425 2.460 0.535 ;
        RECT  2.285 1.200 2.460 1.300 ;
        RECT  2.180 1.200 2.285 1.505 ;
        RECT  1.695 1.395 2.180 1.505 ;
        RECT  2.090 0.315 2.120 0.930 ;
        RECT  2.000 0.315 2.090 1.285 ;
        RECT  1.145 0.315 2.000 0.405 ;
        RECT  0.520 1.180 2.000 1.285 ;
        RECT  0.185 1.395 1.415 1.505 ;
        RECT  0.160 0.390 0.185 0.580 ;
        RECT  0.160 1.195 0.185 1.505 ;
        RECT  0.060 0.390 0.160 1.505 ;
    END
END LHCSNQD2

MACRO LHCSNQD4
    CLASS CORE ;
    FOREIGN LHCSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.370 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.275 4.065 0.695 ;
        RECT  3.955 1.040 4.065 1.490 ;
        RECT  3.850 0.525 3.955 0.695 ;
        RECT  3.850 1.040 3.955 1.210 ;
        RECT  3.550 0.525 3.850 1.210 ;
        RECT  3.435 0.275 3.550 0.695 ;
        RECT  3.435 1.040 3.550 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0802 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.980 1.725 1.090 ;
        RECT  1.150 0.675 1.270 0.775 ;
        RECT  1.050 0.675 1.150 1.090 ;
        RECT  0.350 1.000 1.050 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0415 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.435 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.435 0.585 ;
        RECT  0.650 0.255 0.750 0.585 ;
        RECT  0.480 0.255 0.650 0.365 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.695 ;
        RECT  3.755 -0.165 4.215 0.165 ;
        RECT  3.755 0.325 3.855 0.435 ;
        RECT  3.645 -0.165 3.755 0.435 ;
        RECT  3.285 -0.165 3.645 0.165 ;
        RECT  3.175 -0.165 3.285 0.475 ;
        RECT  2.765 -0.165 3.175 0.165 ;
        RECT  2.655 -0.165 2.765 0.695 ;
        RECT  0.385 -0.165 2.655 0.165 ;
        RECT  0.385 0.475 0.495 0.585 ;
        RECT  0.285 -0.165 0.385 0.585 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.040 4.325 1.965 ;
        RECT  3.805 1.635 4.215 1.965 ;
        RECT  3.695 1.300 3.805 1.965 ;
        RECT  3.285 1.635 3.695 1.965 ;
        RECT  3.175 1.230 3.285 1.965 ;
        RECT  2.765 1.635 3.175 1.965 ;
        RECT  2.655 1.040 2.765 1.965 ;
        RECT  2.630 1.390 2.655 1.965 ;
        RECT  2.385 1.390 2.630 1.500 ;
        RECT  0.000 1.635 2.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.955 0.275 4.065 0.695 ;
        RECT  3.955 1.040 4.065 1.490 ;
        RECT  3.950 0.525 3.955 0.695 ;
        RECT  3.950 1.040 3.955 1.210 ;
        RECT  3.300 0.785 3.440 0.890 ;
        RECT  3.200 0.585 3.300 1.140 ;
        RECT  3.025 0.585 3.200 0.695 ;
        RECT  3.025 1.040 3.200 1.140 ;
        RECT  2.560 0.785 3.075 0.890 ;
        RECT  2.915 0.275 3.025 0.695 ;
        RECT  2.915 1.040 3.025 1.470 ;
        RECT  2.550 0.425 2.560 0.890 ;
        RECT  2.460 0.425 2.550 1.300 ;
        RECT  2.325 0.425 2.460 0.535 ;
        RECT  2.285 1.200 2.460 1.300 ;
        RECT  2.180 1.200 2.285 1.505 ;
        RECT  1.695 1.395 2.180 1.505 ;
        RECT  2.090 0.315 2.120 0.930 ;
        RECT  2.000 0.315 2.090 1.285 ;
        RECT  1.145 0.315 2.000 0.405 ;
        RECT  0.520 1.180 2.000 1.285 ;
        RECT  0.185 1.395 1.415 1.505 ;
        RECT  0.160 0.390 0.185 0.580 ;
        RECT  0.160 1.195 0.185 1.505 ;
        RECT  0.060 0.390 0.160 1.505 ;
    END
END LHCSNQD4

MACRO LHD1
    CLASS CORE ;
    FOREIGN LHD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.275 2.950 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.545 2.555 1.290 ;
        RECT  2.400 0.545 2.445 0.675 ;
        RECT  2.290 1.110 2.445 1.290 ;
        RECT  2.290 0.275 2.400 0.675 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0352 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.710 0.965 1.100 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.885 -0.165 3.000 0.165 ;
        RECT  1.755 -0.165 1.885 0.455 ;
        RECT  0.975 -0.165 1.755 0.165 ;
        RECT  0.805 -0.165 0.975 0.410 ;
        RECT  0.000 -0.165 0.805 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.635 3.000 1.965 ;
        RECT  0.910 1.210 0.985 1.310 ;
        RECT  0.800 1.210 0.910 1.965 ;
        RECT  0.000 1.635 0.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.645 0.730 2.735 1.490 ;
        RECT  2.200 1.400 2.645 1.490 ;
        RECT  2.110 0.275 2.200 1.490 ;
        RECT  2.030 0.275 2.110 0.645 ;
        RECT  2.030 1.245 2.110 1.490 ;
        RECT  1.770 0.545 2.030 0.645 ;
        RECT  1.910 0.755 2.020 1.135 ;
        RECT  1.540 1.045 1.910 1.135 ;
        RECT  1.660 0.545 1.770 0.935 ;
        RECT  1.165 1.435 1.550 1.525 ;
        RECT  1.440 0.275 1.540 1.135 ;
        RECT  1.300 0.275 1.440 0.475 ;
        RECT  1.410 1.045 1.440 1.135 ;
        RECT  1.300 1.045 1.410 1.345 ;
        RECT  1.165 0.585 1.350 0.695 ;
        RECT  1.075 0.500 1.165 1.525 ;
        RECT  0.700 0.500 1.075 0.600 ;
        RECT  0.610 0.500 0.700 1.490 ;
        RECT  0.525 0.500 0.610 0.605 ;
        RECT  0.580 1.210 0.610 1.490 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.365 0.410 1.310 ;
        RECT  0.065 0.365 0.310 0.555 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LHD1

MACRO LHD2
    CLASS CORE ;
    FOREIGN LHD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.150 1.490 ;
        RECT  2.965 0.275 3.050 0.675 ;
        RECT  2.965 1.055 3.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.275 2.585 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0343 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.100 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.635 3.400 1.965 ;
        RECT  0.760 1.335 0.930 1.965 ;
        RECT  0.000 1.635 0.760 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.825 0.790 2.955 0.890 ;
        RECT  2.725 0.790 2.825 1.490 ;
        RECT  2.170 1.400 2.725 1.490 ;
        RECT  2.080 0.275 2.170 1.490 ;
        RECT  1.990 0.275 2.080 0.645 ;
        RECT  1.990 1.245 2.080 1.490 ;
        RECT  1.750 0.545 1.990 0.645 ;
        RECT  1.880 0.755 1.990 1.135 ;
        RECT  1.520 1.045 1.880 1.135 ;
        RECT  1.640 0.545 1.750 0.935 ;
        RECT  1.145 1.435 1.530 1.525 ;
        RECT  1.420 0.275 1.520 1.135 ;
        RECT  1.280 0.275 1.420 0.475 ;
        RECT  1.390 1.045 1.420 1.135 ;
        RECT  1.280 1.045 1.390 1.345 ;
        RECT  1.145 0.585 1.330 0.695 ;
        RECT  1.055 0.365 1.145 1.525 ;
        RECT  0.700 0.365 1.055 0.465 ;
        RECT  0.610 0.365 0.700 1.215 ;
        RECT  0.535 0.365 0.610 0.555 ;
        RECT  0.580 1.025 0.610 1.215 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.365 0.410 1.310 ;
        RECT  0.065 0.365 0.310 0.555 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LHD2

MACRO LHD4
    CLASS CORE ;
    FOREIGN LHD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.310 4.150 0.690 ;
        RECT  4.050 1.110 4.150 1.490 ;
        RECT  3.750 0.310 4.050 1.490 ;
        RECT  3.425 0.310 3.750 0.690 ;
        RECT  3.425 1.110 3.750 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.150 0.690 ;
        RECT  3.050 1.110 3.115 1.290 ;
        RECT  2.750 0.310 3.050 1.290 ;
        RECT  2.425 0.310 2.750 0.690 ;
        RECT  2.425 1.110 2.750 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0343 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.100 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.635 4.400 1.965 ;
        RECT  0.760 1.335 0.930 1.965 ;
        RECT  0.000 1.635 0.760 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.425 0.310 3.650 0.690 ;
        RECT  3.425 1.110 3.650 1.490 ;
        RECT  2.425 0.310 2.650 0.690 ;
        RECT  2.425 1.110 2.650 1.290 ;
        RECT  3.335 0.790 3.550 0.890 ;
        RECT  3.235 0.790 3.335 1.490 ;
        RECT  2.170 1.400 3.235 1.490 ;
        RECT  2.080 0.275 2.170 1.490 ;
        RECT  1.990 0.275 2.080 0.645 ;
        RECT  1.990 1.245 2.080 1.490 ;
        RECT  1.750 0.545 1.990 0.645 ;
        RECT  1.880 0.755 1.990 1.135 ;
        RECT  1.520 1.045 1.880 1.135 ;
        RECT  1.640 0.545 1.750 0.935 ;
        RECT  1.145 1.435 1.530 1.525 ;
        RECT  1.420 0.275 1.520 1.135 ;
        RECT  1.280 0.275 1.420 0.475 ;
        RECT  1.390 1.045 1.420 1.135 ;
        RECT  1.280 1.045 1.390 1.345 ;
        RECT  1.145 0.585 1.330 0.695 ;
        RECT  1.055 0.365 1.145 1.525 ;
        RECT  0.700 0.365 1.055 0.465 ;
        RECT  0.610 0.365 0.700 1.215 ;
        RECT  0.535 0.365 0.610 0.555 ;
        RECT  0.580 1.025 0.610 1.215 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.365 0.410 1.310 ;
        RECT  0.065 0.365 0.310 0.555 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LHD4

MACRO LHQD1
    CLASS CORE ;
    FOREIGN LHQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.275 2.750 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0360 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.965 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.075 -0.165 2.800 0.165 ;
        RECT  0.865 -0.165 1.075 0.405 ;
        RECT  0.510 -0.165 0.865 0.165 ;
        RECT  0.340 -0.165 0.510 0.400 ;
        RECT  0.000 -0.165 0.340 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.975 1.635 2.800 1.965 ;
        RECT  1.865 1.145 1.975 1.965 ;
        RECT  1.085 1.635 1.865 1.965 ;
        RECT  0.975 1.200 1.085 1.965 ;
        RECT  0.875 1.200 0.975 1.310 ;
        RECT  0.510 1.635 0.975 1.965 ;
        RECT  0.340 1.400 0.510 1.965 ;
        RECT  0.000 1.635 0.340 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.290 0.350 2.400 1.295 ;
        RECT  2.070 0.725 2.180 1.055 ;
        RECT  1.630 0.965 2.070 1.055 ;
        RECT  1.770 0.350 1.880 0.875 ;
        RECT  1.430 1.435 1.640 1.545 ;
        RECT  1.540 0.310 1.630 1.055 ;
        RECT  1.415 0.310 1.540 0.500 ;
        RECT  1.525 0.965 1.540 1.055 ;
        RECT  1.415 0.965 1.525 1.325 ;
        RECT  1.325 0.610 1.450 0.710 ;
        RECT  1.325 1.435 1.430 1.525 ;
        RECT  1.215 0.495 1.325 1.525 ;
        RECT  0.760 0.495 1.215 0.600 ;
        RECT  0.655 0.495 0.760 1.470 ;
        RECT  0.430 0.490 0.540 1.310 ;
        RECT  0.055 0.490 0.430 0.600 ;
        RECT  0.195 1.200 0.430 1.310 ;
        RECT  0.085 1.200 0.195 1.460 ;
        RECT  1.880 0.350 2.290 0.460 ;
        RECT  2.085 1.185 2.290 1.295 ;
    END
END LHQD1

MACRO LHQD2
    CLASS CORE ;
    FOREIGN LHQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.275 2.750 1.490 ;
        RECT  2.565 0.275 2.650 0.695 ;
        RECT  2.565 1.040 2.650 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0367 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.965 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.635 3.000 1.965 ;
        RECT  1.830 1.145 1.940 1.965 ;
        RECT  0.995 1.635 1.830 1.965 ;
        RECT  0.825 1.345 0.995 1.965 ;
        RECT  0.000 1.635 0.825 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.255 0.350 2.365 1.295 ;
        RECT  1.845 0.350 2.255 0.460 ;
        RECT  2.050 1.185 2.255 1.295 ;
        RECT  2.035 0.725 2.145 1.055 ;
        RECT  1.595 0.965 2.035 1.055 ;
        RECT  1.735 0.350 1.845 0.875 ;
        RECT  1.395 1.435 1.605 1.545 ;
        RECT  1.505 0.310 1.595 1.055 ;
        RECT  1.380 0.310 1.505 0.500 ;
        RECT  1.490 0.965 1.505 1.055 ;
        RECT  1.380 0.965 1.490 1.325 ;
        RECT  1.290 0.610 1.415 0.710 ;
        RECT  1.290 1.435 1.395 1.525 ;
        RECT  1.180 0.275 1.290 1.525 ;
        RECT  0.745 0.275 1.180 0.380 ;
        RECT  0.650 0.275 0.745 1.215 ;
        RECT  0.430 0.500 0.540 1.300 ;
        RECT  0.055 0.500 0.430 0.600 ;
        RECT  0.195 1.200 0.430 1.300 ;
        RECT  0.085 1.200 0.195 1.450 ;
    END
END LHQD2

MACRO LHQD4
    CLASS CORE ;
    FOREIGN LHQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.150 0.690 ;
        RECT  3.050 1.110 3.150 1.490 ;
        RECT  2.750 0.310 3.050 1.490 ;
        RECT  2.425 0.310 2.750 0.690 ;
        RECT  2.425 1.110 2.750 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0343 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.100 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.165 3.400 0.165 ;
        RECT  0.760 -0.165 0.930 0.285 ;
        RECT  0.000 -0.165 0.760 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.635 3.400 1.965 ;
        RECT  0.760 1.335 0.930 1.965 ;
        RECT  0.000 1.635 0.760 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.425 0.310 2.650 0.690 ;
        RECT  2.425 1.110 2.650 1.490 ;
        RECT  2.080 0.310 2.170 1.295 ;
        RECT  1.750 0.310 2.080 0.410 ;
        RECT  1.945 1.185 2.080 1.295 ;
        RECT  1.880 0.755 1.990 1.085 ;
        RECT  1.520 0.995 1.880 1.085 ;
        RECT  1.640 0.310 1.750 0.905 ;
        RECT  1.145 1.435 1.530 1.525 ;
        RECT  1.420 0.275 1.520 1.085 ;
        RECT  1.280 0.275 1.420 0.475 ;
        RECT  1.390 0.995 1.420 1.085 ;
        RECT  1.280 0.995 1.390 1.345 ;
        RECT  1.145 0.585 1.330 0.695 ;
        RECT  1.055 0.375 1.145 1.525 ;
        RECT  0.700 0.375 1.055 0.475 ;
        RECT  0.610 0.375 0.700 1.215 ;
        RECT  0.535 0.375 0.610 0.575 ;
        RECT  0.580 1.025 0.610 1.215 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.365 0.410 1.310 ;
        RECT  0.065 0.365 0.310 0.555 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LHQD4

MACRO LHSND1
    CLASS CORE ;
    FOREIGN LHSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.770 1.100 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.500 2.650 0.690 ;
        RECT  2.550 1.025 2.645 1.125 ;
        RECT  2.450 0.500 2.550 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.285 3.150 1.490 ;
        RECT  3.025 0.285 3.050 0.675 ;
        RECT  3.025 0.995 3.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0491 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.000 1.080 1.105 ;
        RECT  0.675 0.525 0.780 1.105 ;
        RECT  0.350 1.000 0.675 1.105 ;
        RECT  0.240 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.500 0.565 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.870 -0.165 3.200 0.165 ;
        RECT  2.760 -0.165 2.870 0.645 ;
        RECT  2.110 -0.165 2.760 0.165 ;
        RECT  1.960 -0.165 2.110 0.345 ;
        RECT  1.390 -0.165 1.960 0.165 ;
        RECT  1.280 -0.165 1.390 0.660 ;
        RECT  0.000 -0.165 1.280 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.635 3.200 1.965 ;
        RECT  2.715 1.395 2.905 1.965 ;
        RECT  2.035 1.635 2.715 1.965 ;
        RECT  1.865 1.420 2.035 1.965 ;
        RECT  0.000 1.635 1.865 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.860 0.755 2.940 0.925 ;
        RECT  2.760 0.755 2.860 1.305 ;
        RECT  2.325 1.215 2.760 1.305 ;
        RECT  2.325 0.310 2.415 0.410 ;
        RECT  2.225 0.310 2.325 1.490 ;
        RECT  2.015 0.460 2.115 1.310 ;
        RECT  1.715 0.460 2.015 0.560 ;
        RECT  1.690 1.210 2.015 1.310 ;
        RECT  1.570 1.210 1.690 1.525 ;
        RECT  1.090 1.425 1.570 1.525 ;
        RECT  1.325 0.750 1.520 0.920 ;
        RECT  1.235 0.750 1.325 1.295 ;
        RECT  1.115 0.750 1.235 0.840 ;
        RECT  0.725 1.205 1.235 1.295 ;
        RECT  1.025 0.295 1.115 0.840 ;
        RECT  0.735 0.295 1.025 0.425 ;
        RECT  0.175 1.425 0.840 1.525 ;
        RECT  0.150 0.275 0.195 0.510 ;
        RECT  0.150 1.200 0.175 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LHSND1

MACRO LHSND2
    CLASS CORE ;
    FOREIGN LHSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0415 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.605 1.760 1.100 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.265 2.785 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.275 3.350 1.515 ;
        RECT  3.160 0.275 3.250 0.655 ;
        RECT  3.160 1.040 3.250 1.515 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0491 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.000 1.080 1.105 ;
        RECT  0.675 0.525 0.790 1.105 ;
        RECT  0.350 1.000 0.675 1.105 ;
        RECT  0.240 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.500 0.565 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.375 -0.165 3.600 0.165 ;
        RECT  1.245 -0.165 1.375 0.465 ;
        RECT  0.000 -0.165 1.245 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.045 1.635 3.600 1.965 ;
        RECT  2.875 1.395 3.045 1.965 ;
        RECT  1.985 1.635 2.875 1.965 ;
        RECT  1.815 1.420 1.985 1.965 ;
        RECT  0.000 1.635 1.815 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.040 0.780 3.160 0.890 ;
        RECT  2.930 0.780 3.040 1.305 ;
        RECT  2.300 1.215 2.930 1.305 ;
        RECT  2.150 0.260 2.300 1.490 ;
        RECT  1.905 0.350 2.015 1.310 ;
        RECT  1.665 0.350 1.905 0.450 ;
        RECT  1.660 1.210 1.905 1.310 ;
        RECT  1.540 1.210 1.660 1.525 ;
        RECT  1.090 1.425 1.540 1.525 ;
        RECT  1.325 0.905 1.500 1.075 ;
        RECT  1.235 0.575 1.325 1.295 ;
        RECT  1.125 0.575 1.235 0.665 ;
        RECT  0.725 1.205 1.235 1.295 ;
        RECT  1.035 0.295 1.125 0.665 ;
        RECT  0.735 0.295 1.035 0.425 ;
        RECT  0.175 1.425 0.840 1.525 ;
        RECT  0.140 0.275 0.195 0.510 ;
        RECT  0.140 1.200 0.175 1.525 ;
        RECT  0.050 0.275 0.140 1.525 ;
    END
END LHSND2

MACRO LHSND4
    CLASS CORE ;
    FOREIGN LHSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.700 1.950 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.310 3.695 0.695 ;
        RECT  3.450 1.110 3.695 1.290 ;
        RECT  3.150 0.310 3.450 1.290 ;
        RECT  3.005 0.310 3.150 0.695 ;
        RECT  3.005 1.110 3.150 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.310 4.695 0.690 ;
        RECT  4.650 1.110 4.695 1.490 ;
        RECT  4.350 0.310 4.650 1.490 ;
        RECT  4.005 0.310 4.350 0.690 ;
        RECT  4.005 1.110 4.350 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0765 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.000 1.150 1.105 ;
        RECT  0.730 0.510 0.840 1.105 ;
        RECT  0.350 1.000 0.730 1.105 ;
        RECT  0.240 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.580 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.915 -0.165 5.000 0.165 ;
        RECT  4.805 -0.165 4.915 0.690 ;
        RECT  0.500 -0.165 4.805 0.165 ;
        RECT  0.310 -0.165 0.500 0.415 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.915 1.635 5.000 1.965 ;
        RECT  4.805 1.110 4.915 1.965 ;
        RECT  0.000 1.635 4.805 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.005 0.310 4.250 0.690 ;
        RECT  4.005 1.110 4.250 1.490 ;
        RECT  3.550 0.310 3.695 0.695 ;
        RECT  3.550 1.110 3.695 1.290 ;
        RECT  3.005 0.310 3.050 0.695 ;
        RECT  3.005 1.110 3.050 1.290 ;
        RECT  3.895 0.800 4.140 0.910 ;
        RECT  3.805 0.800 3.895 1.505 ;
        RECT  2.655 1.400 3.805 1.505 ;
        RECT  2.760 0.600 2.870 1.200 ;
        RECT  2.655 0.600 2.760 0.690 ;
        RECT  2.655 1.110 2.760 1.200 ;
        RECT  2.545 0.310 2.655 0.690 ;
        RECT  2.545 1.110 2.655 1.505 ;
        RECT  2.455 0.800 2.650 0.910 ;
        RECT  2.345 0.345 2.455 1.505 ;
        RECT  1.745 0.345 2.345 0.455 ;
        RECT  1.695 1.395 2.345 1.505 ;
        RECT  2.125 0.700 2.235 1.295 ;
        RECT  1.500 1.205 2.125 1.295 ;
        RECT  1.505 1.395 1.695 1.525 ;
        RECT  1.090 1.425 1.505 1.525 ;
        RECT  1.390 0.305 1.500 1.295 ;
        RECT  0.780 0.305 1.390 0.415 ;
        RECT  0.725 1.205 1.390 1.295 ;
        RECT  0.175 1.425 0.840 1.525 ;
        RECT  0.140 0.275 0.195 0.510 ;
        RECT  0.140 1.200 0.175 1.525 ;
        RECT  0.050 0.275 0.140 1.525 ;
    END
END LHSND4

MACRO LHSNDD1
    CLASS CORE ;
    FOREIGN LHSNDD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.170 0.710 2.250 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.305 3.150 1.175 ;
        RECT  2.865 0.305 3.050 0.415 ;
        RECT  2.915 0.965 3.050 1.175 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.275 3.550 1.490 ;
        RECT  3.415 0.275 3.450 0.675 ;
        RECT  3.420 1.080 3.450 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.600 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.635 3.600 1.965 ;
        RECT  2.350 1.495 2.520 1.965 ;
        RECT  0.000 1.635 2.350 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.330 0.750 3.360 0.920 ;
        RECT  3.240 0.750 3.330 1.375 ;
        RECT  2.810 1.285 3.240 1.375 ;
        RECT  2.700 0.495 2.810 1.460 ;
        RECT  2.480 0.500 2.590 1.300 ;
        RECT  2.205 0.500 2.480 0.610 ;
        RECT  2.185 1.200 2.480 1.300 ;
        RECT  2.075 1.200 2.185 1.525 ;
        RECT  1.620 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.020 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.265 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.625 1.115 ;
        RECT  1.155 1.435 1.365 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.700 1.020 1.190 1.115 ;
        RECT  0.460 1.435 1.155 1.525 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHSNDD1

MACRO LHSNDD2
    CLASS CORE ;
    FOREIGN LHSNDD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.710 2.350 1.090 ;
        RECT  2.170 0.710 2.240 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.175 1.250 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.275 3.750 1.490 ;
        RECT  3.565 0.275 3.650 0.675 ;
        RECT  3.565 1.080 3.650 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 4.000 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.420 0.780 3.560 0.890 ;
        RECT  3.330 0.780 3.420 1.480 ;
        RECT  2.940 1.370 3.330 1.480 ;
        RECT  2.840 0.305 2.940 1.480 ;
        RECT  2.515 0.305 2.840 0.415 ;
        RECT  2.515 1.370 2.840 1.480 ;
        RECT  2.620 0.510 2.730 1.280 ;
        RECT  2.265 0.510 2.620 0.620 ;
        RECT  2.185 1.180 2.620 1.280 ;
        RECT  2.075 1.180 2.185 1.525 ;
        RECT  1.620 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.030 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.265 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.625 1.115 ;
        RECT  1.155 1.435 1.365 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.700 1.020 1.190 1.115 ;
        RECT  0.460 1.435 1.155 1.525 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHSNDD2

MACRO LHSNDD4
    CLASS CORE ;
    FOREIGN LHSNDD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.700 2.360 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.325 4.265 0.635 ;
        RECT  4.050 1.110 4.255 1.290 ;
        RECT  3.750 0.325 4.050 1.290 ;
        RECT  3.545 0.325 3.750 0.635 ;
        RECT  3.555 1.110 3.750 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.230 0.325 5.285 0.635 ;
        RECT  5.230 1.100 5.285 1.410 ;
        RECT  4.930 0.325 5.230 1.410 ;
        RECT  4.565 0.325 4.930 0.635 ;
        RECT  4.565 1.100 4.930 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.495 -0.165 5.600 0.165 ;
        RECT  5.385 -0.165 5.495 0.685 ;
        RECT  0.000 -0.165 5.385 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.495 1.635 5.600 1.965 ;
        RECT  5.385 1.050 5.495 1.965 ;
        RECT  0.000 1.635 5.385 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.565 0.325 4.850 0.635 ;
        RECT  4.565 1.100 4.850 1.410 ;
        RECT  4.150 0.325 4.265 0.635 ;
        RECT  4.150 1.110 4.255 1.290 ;
        RECT  3.545 0.325 3.650 0.635 ;
        RECT  3.555 1.110 3.650 1.290 ;
        RECT  4.465 0.780 4.710 0.890 ;
        RECT  4.375 0.780 4.465 1.505 ;
        RECT  3.195 1.400 4.375 1.505 ;
        RECT  3.310 0.595 3.410 1.150 ;
        RECT  3.195 0.595 3.310 0.685 ;
        RECT  3.195 1.050 3.310 1.150 ;
        RECT  3.085 0.275 3.195 0.685 ;
        RECT  3.085 1.050 3.195 1.505 ;
        RECT  2.995 0.780 3.190 0.890 ;
        RECT  2.885 0.490 2.995 1.495 ;
        RECT  2.275 0.490 2.885 0.600 ;
        RECT  1.830 1.385 2.885 1.495 ;
        RECT  2.660 0.750 2.770 1.295 ;
        RECT  2.030 1.205 2.660 1.295 ;
        RECT  1.920 0.295 2.030 1.295 ;
        RECT  1.235 0.295 1.920 0.405 ;
        RECT  1.475 1.205 1.920 1.295 ;
        RECT  1.620 1.385 1.830 1.525 ;
        RECT  1.300 1.005 1.625 1.115 ;
        RECT  1.265 1.205 1.475 1.315 ;
        RECT  1.155 1.435 1.365 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.700 1.020 1.190 1.115 ;
        RECT  0.460 1.435 1.155 1.525 ;
        RECT  0.610 0.275 0.700 1.240 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.030 0.610 1.240 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHSNDD4

MACRO LHSNDQD1
    CLASS CORE ;
    FOREIGN LHSNDQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.170 0.710 2.250 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.150 1.490 ;
        RECT  3.015 0.275 3.050 0.675 ;
        RECT  3.015 1.080 3.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.200 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.200 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 0.750 2.960 0.920 ;
        RECT  2.820 0.305 2.920 1.495 ;
        RECT  2.465 0.305 2.820 0.415 ;
        RECT  2.485 1.385 2.820 1.495 ;
        RECT  2.600 0.510 2.710 1.290 ;
        RECT  2.215 0.510 2.600 0.620 ;
        RECT  2.165 1.190 2.600 1.290 ;
        RECT  2.055 1.190 2.165 1.525 ;
        RECT  1.600 1.415 2.055 1.525 ;
        RECT  1.920 0.750 2.010 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.245 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.605 1.115 ;
        RECT  1.135 1.435 1.345 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.700 1.020 1.190 1.115 ;
        RECT  0.460 1.435 1.135 1.525 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHSNDQD1

MACRO LHSNDQD2
    CLASS CORE ;
    FOREIGN LHSNDQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.220 0.710 2.250 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.575 3.350 1.180 ;
        RECT  3.205 0.575 3.250 0.675 ;
        RECT  3.205 1.080 3.250 1.180 ;
        RECT  3.095 0.275 3.205 0.675 ;
        RECT  3.095 1.080 3.205 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 -0.165 3.600 0.165 ;
        RECT  3.355 -0.165 3.465 0.485 ;
        RECT  0.880 -0.165 3.355 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 1.635 3.600 1.965 ;
        RECT  3.355 1.280 3.465 1.965 ;
        RECT  0.000 1.635 3.355 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.000 0.780 3.160 0.890 ;
        RECT  2.900 0.305 3.000 1.495 ;
        RECT  2.525 0.305 2.900 0.415 ;
        RECT  2.545 1.385 2.900 1.495 ;
        RECT  2.660 0.510 2.770 1.290 ;
        RECT  2.275 0.510 2.660 0.620 ;
        RECT  2.185 1.190 2.660 1.290 ;
        RECT  2.075 1.190 2.185 1.525 ;
        RECT  1.600 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.020 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.245 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.605 1.115 ;
        RECT  1.135 1.435 1.345 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.700 1.020 1.190 1.115 ;
        RECT  0.460 1.435 1.135 1.525 ;
        RECT  0.610 0.440 0.700 1.340 ;
        RECT  0.575 0.440 0.610 0.650 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHSNDQD2

MACRO LHSNDQD4
    CLASS CORE ;
    FOREIGN LHSNDQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.220 0.710 2.250 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.325 3.750 0.635 ;
        RECT  3.650 1.100 3.750 1.410 ;
        RECT  3.350 0.325 3.650 1.410 ;
        RECT  3.015 0.325 3.350 0.635 ;
        RECT  3.015 1.100 3.350 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.280 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.015 0.325 3.250 0.635 ;
        RECT  3.015 1.100 3.250 1.410 ;
        RECT  2.905 0.780 3.160 0.890 ;
        RECT  2.805 0.305 2.905 1.495 ;
        RECT  2.515 0.305 2.805 0.415 ;
        RECT  2.535 1.385 2.805 1.495 ;
        RECT  2.585 0.510 2.695 1.290 ;
        RECT  2.265 0.510 2.585 0.620 ;
        RECT  2.185 1.190 2.585 1.290 ;
        RECT  2.075 1.190 2.185 1.525 ;
        RECT  1.600 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.020 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.245 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.605 1.115 ;
        RECT  1.135 1.435 1.345 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.700 1.020 1.190 1.115 ;
        RECT  0.460 1.435 1.135 1.525 ;
        RECT  0.610 0.275 0.700 1.340 ;
        RECT  0.575 0.275 0.610 0.675 ;
        RECT  0.575 1.130 0.610 1.340 ;
        RECT  0.460 0.750 0.520 0.920 ;
        RECT  0.370 0.490 0.460 1.525 ;
        RECT  0.045 0.490 0.370 0.600 ;
        RECT  0.045 1.200 0.370 1.310 ;
    END
END LHSNDQD4

MACRO LHSNQD1
    CLASS CORE ;
    FOREIGN LHSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.770 1.100 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.785 0.285 2.950 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0491 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.000 1.080 1.105 ;
        RECT  0.680 0.525 0.790 1.105 ;
        RECT  0.350 1.000 0.680 1.105 ;
        RECT  0.240 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.500 0.565 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.650 -0.165 3.000 0.165 ;
        RECT  2.510 -0.165 2.650 0.645 ;
        RECT  2.130 -0.165 2.510 0.165 ;
        RECT  1.940 -0.165 2.130 0.335 ;
        RECT  1.400 -0.165 1.940 0.165 ;
        RECT  1.270 -0.165 1.400 0.660 ;
        RECT  0.000 -0.165 1.270 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.645 1.635 3.000 1.965 ;
        RECT  2.510 1.040 2.645 1.965 ;
        RECT  2.035 1.635 2.510 1.965 ;
        RECT  1.865 1.420 2.035 1.965 ;
        RECT  0.000 1.635 1.865 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.375 0.740 2.675 0.930 ;
        RECT  2.340 0.275 2.375 0.930 ;
        RECT  2.225 0.275 2.340 1.490 ;
        RECT  1.980 0.445 2.100 1.310 ;
        RECT  1.715 0.445 1.980 0.575 ;
        RECT  1.700 1.210 1.980 1.310 ;
        RECT  1.580 1.210 1.700 1.525 ;
        RECT  1.090 1.425 1.580 1.525 ;
        RECT  1.325 0.750 1.520 0.920 ;
        RECT  1.235 0.750 1.325 1.295 ;
        RECT  1.115 0.750 1.235 0.840 ;
        RECT  0.725 1.205 1.235 1.295 ;
        RECT  1.025 0.295 1.115 0.840 ;
        RECT  0.735 0.295 1.025 0.425 ;
        RECT  0.175 1.425 0.840 1.525 ;
        RECT  0.150 0.275 0.195 0.510 ;
        RECT  0.150 1.200 0.175 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LHSNQD1

MACRO LHSNQD2
    CLASS CORE ;
    FOREIGN LHSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.770 1.100 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.875 0.545 2.950 1.155 ;
        RECT  2.850 0.265 2.875 1.515 ;
        RECT  2.745 0.265 2.850 0.695 ;
        RECT  2.745 1.035 2.850 1.515 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0491 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.000 1.080 1.105 ;
        RECT  0.680 0.525 0.790 1.105 ;
        RECT  0.350 1.000 0.680 1.105 ;
        RECT  0.240 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.500 0.565 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.135 -0.165 3.200 0.165 ;
        RECT  3.005 -0.165 3.135 0.445 ;
        RECT  2.615 -0.165 3.005 0.165 ;
        RECT  2.495 -0.165 2.615 0.695 ;
        RECT  2.100 -0.165 2.495 0.165 ;
        RECT  1.970 -0.165 2.100 0.345 ;
        RECT  1.390 -0.165 1.970 0.165 ;
        RECT  1.280 -0.165 1.390 0.660 ;
        RECT  0.000 -0.165 1.280 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.135 1.635 3.200 1.965 ;
        RECT  3.005 1.275 3.135 1.965 ;
        RECT  2.615 1.635 3.005 1.965 ;
        RECT  2.485 1.035 2.615 1.965 ;
        RECT  2.035 1.635 2.485 1.965 ;
        RECT  1.865 1.420 2.035 1.965 ;
        RECT  0.000 1.635 1.865 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.335 0.810 2.740 0.925 ;
        RECT  2.335 0.310 2.405 0.410 ;
        RECT  2.215 0.310 2.335 1.490 ;
        RECT  1.990 0.460 2.100 1.310 ;
        RECT  1.715 0.460 1.990 0.560 ;
        RECT  1.690 1.210 1.990 1.310 ;
        RECT  1.570 1.210 1.690 1.525 ;
        RECT  1.090 1.425 1.570 1.525 ;
        RECT  1.325 0.750 1.520 0.920 ;
        RECT  1.115 0.750 1.235 0.840 ;
        RECT  0.725 1.205 1.235 1.295 ;
        RECT  1.025 0.295 1.115 0.840 ;
        RECT  0.735 0.295 1.025 0.425 ;
        RECT  0.175 1.425 0.840 1.525 ;
        RECT  0.150 0.275 0.195 0.510 ;
        RECT  0.150 1.200 0.175 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
        RECT  1.235 0.750 1.325 1.295 ;
    END
END LHSNQD2

MACRO LHSNQD4
    CLASS CORE ;
    FOREIGN LHSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.510 1.950 0.920 ;
        RECT  1.760 0.730 1.845 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.505 3.270 0.675 ;
        RECT  3.110 0.990 3.240 1.515 ;
        RECT  3.050 0.990 3.110 1.160 ;
        RECT  2.750 0.505 3.050 1.160 ;
        RECT  2.550 0.505 2.750 0.675 ;
        RECT  2.720 0.990 2.750 1.160 ;
        RECT  2.590 0.990 2.720 1.515 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0765 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.000 1.100 1.105 ;
        RECT  0.730 0.510 0.840 1.105 ;
        RECT  0.350 1.000 0.730 1.105 ;
        RECT  0.240 0.710 0.350 1.105 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.580 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 -0.165 3.600 0.165 ;
        RECT  0.310 -0.165 0.500 0.415 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.490 1.635 3.600 1.965 ;
        RECT  3.380 1.055 3.490 1.965 ;
        RECT  2.980 1.635 3.380 1.965 ;
        RECT  2.850 1.270 2.980 1.965 ;
        RECT  2.480 1.635 2.850 1.965 ;
        RECT  2.295 1.390 2.480 1.965 ;
        RECT  1.970 1.635 2.295 1.965 ;
        RECT  1.800 1.405 1.970 1.965 ;
        RECT  0.000 1.635 1.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 0.505 3.270 0.675 ;
        RECT  3.150 0.990 3.240 1.515 ;
        RECT  2.550 0.505 2.650 0.675 ;
        RECT  2.590 0.990 2.650 1.515 ;
        RECT  3.400 0.275 3.520 0.890 ;
        RECT  2.165 0.275 3.400 0.380 ;
        RECT  3.255 0.765 3.400 0.890 ;
        RECT  2.315 0.750 2.420 1.295 ;
        RECT  2.260 0.750 2.315 0.920 ;
        RECT  1.670 1.205 2.315 1.295 ;
        RECT  2.165 1.025 2.205 1.115 ;
        RECT  2.060 0.275 2.165 1.115 ;
        RECT  2.035 1.025 2.060 1.115 ;
        RECT  1.670 0.330 1.915 0.420 ;
        RECT  1.580 0.330 1.670 1.525 ;
        RECT  1.540 1.045 1.580 1.525 ;
        RECT  1.090 1.425 1.540 1.525 ;
        RECT  1.340 0.750 1.490 0.920 ;
        RECT  1.230 0.305 1.340 1.295 ;
        RECT  0.780 0.305 1.230 0.415 ;
        RECT  0.175 1.425 0.840 1.525 ;
        RECT  0.140 0.275 0.195 0.510 ;
        RECT  0.140 1.200 0.175 1.525 ;
        RECT  0.050 0.275 0.140 1.525 ;
        RECT  0.725 1.205 1.230 1.295 ;
    END
END LHSNQD4

MACRO LNCND1
    CLASS CORE ;
    FOREIGN LNCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1330 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.025 3.065 1.125 ;
        RECT  2.950 0.480 3.055 0.650 ;
        RECT  2.850 0.480 2.950 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.425 0.285 3.550 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.495 ;
        RECT  1.110 1.345 1.200 1.495 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.710 0.355 1.435 ;
        RECT  0.245 0.710 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 -0.165 3.600 0.165 ;
        RECT  3.100 -0.165 3.270 0.285 ;
        RECT  2.760 -0.165 3.100 0.165 ;
        RECT  2.660 -0.165 2.760 0.685 ;
        RECT  0.000 -0.165 2.660 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.635 3.600 1.965 ;
        RECT  3.100 1.415 3.270 1.965 ;
        RECT  2.805 1.635 3.100 1.965 ;
        RECT  2.615 1.395 2.805 1.965 ;
        RECT  0.000 1.635 2.615 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.180 0.730 3.295 1.305 ;
        RECT  2.570 1.215 3.180 1.305 ;
        RECT  2.500 0.305 2.570 1.305 ;
        RECT  2.470 0.305 2.500 1.465 ;
        RECT  2.355 0.305 2.470 0.405 ;
        RECT  2.400 1.215 2.470 1.465 ;
        RECT  2.290 0.740 2.380 0.930 ;
        RECT  2.190 0.495 2.290 1.495 ;
        RECT  1.680 1.395 2.190 1.495 ;
        RECT  2.000 0.315 2.100 1.255 ;
        RECT  1.135 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.710 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.600 ;
        RECT  0.155 0.405 0.210 0.600 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.405 0.155 1.515 ;
    END
END LNCND1

MACRO LNCND2
    CLASS CORE ;
    FOREIGN LNCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.275 2.975 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.465 0.510 3.550 1.195 ;
        RECT  3.450 0.275 3.465 1.490 ;
        RECT  3.355 0.275 3.450 0.675 ;
        RECT  3.355 1.045 3.450 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.425 1.415 1.400 1.525 ;
        RECT  0.355 1.175 0.425 1.525 ;
        RECT  0.335 0.710 0.355 1.525 ;
        RECT  0.240 0.710 0.335 1.265 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0406 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.495 1.875 0.665 ;
        RECT  1.445 0.495 1.555 0.890 ;
        RECT  0.750 0.495 1.445 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.445 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.165 3.800 0.165 ;
        RECT  3.615 -0.165 3.725 0.445 ;
        RECT  0.000 -0.165 3.615 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.635 3.800 1.965 ;
        RECT  3.610 1.325 3.730 1.965 ;
        RECT  0.000 1.635 3.610 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.210 0.785 3.360 0.885 ;
        RECT  3.120 0.785 3.210 1.505 ;
        RECT  2.555 1.395 3.120 1.505 ;
        RECT  2.455 0.305 2.555 1.505 ;
        RECT  2.300 0.305 2.455 0.415 ;
        RECT  2.365 1.315 2.455 1.505 ;
        RECT  2.255 0.505 2.340 1.215 ;
        RECT  2.240 0.505 2.255 1.525 ;
        RECT  2.145 0.505 2.240 0.685 ;
        RECT  2.145 1.035 2.240 1.525 ;
        RECT  1.660 1.415 2.145 1.525 ;
        RECT  2.055 0.775 2.100 0.945 ;
        RECT  1.965 0.315 2.055 1.305 ;
        RECT  1.115 0.315 1.965 0.405 ;
        RECT  0.515 1.195 1.965 1.305 ;
        RECT  1.355 1.000 1.690 1.105 ;
        RECT  1.245 0.675 1.355 1.105 ;
        RECT  1.040 0.675 1.245 0.785 ;
        RECT  0.555 0.985 1.245 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.205 0.495 0.445 0.600 ;
        RECT  0.150 1.355 0.225 1.525 ;
        RECT  0.150 0.405 0.205 0.600 ;
        RECT  0.060 0.405 0.150 1.525 ;
    END
END LNCND2

MACRO LNCND4
    CLASS CORE ;
    FOREIGN LNCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.310 3.845 0.690 ;
        RECT  3.650 1.110 3.845 1.290 ;
        RECT  3.350 0.310 3.650 1.290 ;
        RECT  3.135 0.310 3.350 0.690 ;
        RECT  3.135 1.110 3.350 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.310 4.885 0.690 ;
        RECT  4.850 1.110 4.885 1.490 ;
        RECT  4.550 0.310 4.850 1.490 ;
        RECT  4.175 0.310 4.550 0.690 ;
        RECT  4.175 1.110 4.550 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0812 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.425 1.415 1.390 1.525 ;
        RECT  0.355 1.175 0.425 1.525 ;
        RECT  0.335 0.700 0.355 1.525 ;
        RECT  0.240 0.700 0.335 1.265 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0406 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.495 1.875 0.665 ;
        RECT  1.445 0.495 1.555 0.890 ;
        RECT  0.750 0.495 1.445 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.445 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 -0.165 5.200 0.165 ;
        RECT  4.995 -0.165 5.105 0.690 ;
        RECT  4.065 -0.165 4.995 0.165 ;
        RECT  3.955 -0.165 4.065 0.690 ;
        RECT  3.025 -0.165 3.955 0.165 ;
        RECT  2.915 -0.165 3.025 0.465 ;
        RECT  2.505 -0.165 2.915 0.165 ;
        RECT  2.395 -0.165 2.505 0.465 ;
        RECT  0.000 -0.165 2.395 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 1.635 5.200 1.965 ;
        RECT  4.995 1.110 5.105 1.965 ;
        RECT  2.505 1.635 4.995 1.965 ;
        RECT  2.395 1.305 2.505 1.965 ;
        RECT  0.000 1.635 2.395 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.175 0.310 4.450 0.690 ;
        RECT  4.175 1.110 4.450 1.490 ;
        RECT  3.750 0.310 3.845 0.690 ;
        RECT  3.750 1.110 3.845 1.290 ;
        RECT  3.135 0.310 3.250 0.690 ;
        RECT  3.135 1.110 3.250 1.290 ;
        RECT  4.065 0.800 4.320 0.900 ;
        RECT  3.955 0.800 4.065 1.525 ;
        RECT  2.875 1.415 3.955 1.525 ;
        RECT  2.765 0.555 2.875 1.525 ;
        RECT  2.655 0.310 2.765 0.690 ;
        RECT  2.655 1.110 2.765 1.525 ;
        RECT  2.340 0.800 2.660 0.900 ;
        RECT  2.255 0.555 2.340 1.210 ;
        RECT  2.240 0.310 2.255 1.525 ;
        RECT  2.145 0.310 2.240 0.685 ;
        RECT  2.145 1.110 2.240 1.525 ;
        RECT  1.670 1.415 2.145 1.525 ;
        RECT  2.055 0.775 2.100 0.945 ;
        RECT  1.965 0.315 2.055 1.305 ;
        RECT  1.125 0.315 1.965 0.405 ;
        RECT  0.515 1.195 1.965 1.305 ;
        RECT  1.355 1.000 1.680 1.105 ;
        RECT  1.245 0.675 1.355 1.105 ;
        RECT  1.040 0.675 1.245 0.785 ;
        RECT  0.555 0.985 1.245 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.205 0.495 0.445 0.585 ;
        RECT  0.150 1.355 0.225 1.525 ;
        RECT  0.150 0.390 0.205 0.585 ;
        RECT  0.060 0.390 0.150 1.525 ;
    END
END LNCND4

MACRO LNCNDD1
    CLASS CORE ;
    FOREIGN LNCNDD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1210 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.525 3.310 0.635 ;
        RECT  3.150 1.020 3.310 1.130 ;
        RECT  3.050 0.525 3.150 1.130 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.275 3.750 1.490 ;
        RECT  3.615 0.275 3.650 0.685 ;
        RECT  3.615 1.080 3.650 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.800 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.415 0.305 3.525 1.340 ;
        RECT  2.610 0.305 3.415 0.415 ;
        RECT  2.770 1.240 3.415 1.340 ;
        RECT  2.585 0.780 2.940 0.890 ;
        RECT  2.660 1.240 2.770 1.525 ;
        RECT  2.565 0.505 2.585 0.890 ;
        RECT  2.475 0.505 2.565 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.280 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.280 0.405 ;
        RECT  0.795 1.205 2.280 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCNDD1

MACRO LNCNDD2
    CLASS CORE ;
    FOREIGN LNCNDD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.525 3.350 1.130 ;
        RECT  3.150 0.525 3.250 0.635 ;
        RECT  3.150 1.020 3.250 1.130 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.585 3.950 1.180 ;
        RECT  3.830 0.585 3.850 0.685 ;
        RECT  3.830 1.080 3.850 1.180 ;
        RECT  3.720 0.275 3.830 0.685 ;
        RECT  3.720 1.080 3.830 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0419 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.090 -0.165 4.200 0.165 ;
        RECT  3.980 -0.165 4.090 0.485 ;
        RECT  0.880 -0.165 3.980 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.090 1.635 4.200 1.965 ;
        RECT  3.980 1.280 4.090 1.965 ;
        RECT  3.600 1.635 3.980 1.965 ;
        RECT  3.430 1.400 3.600 1.965 ;
        RECT  3.080 1.635 3.430 1.965 ;
        RECT  2.910 1.400 3.080 1.965 ;
        RECT  0.000 1.635 2.910 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.630 0.780 3.755 0.890 ;
        RECT  3.520 0.305 3.630 1.310 ;
        RECT  2.640 0.305 3.520 0.415 ;
        RECT  2.800 1.220 3.520 1.310 ;
        RECT  2.615 0.780 3.060 0.890 ;
        RECT  2.690 1.220 2.800 1.525 ;
        RECT  2.595 0.505 2.615 0.890 ;
        RECT  2.505 0.505 2.595 1.525 ;
        RECT  2.010 1.415 2.505 1.525 ;
        RECT  2.320 0.295 2.410 1.315 ;
        RECT  1.465 0.295 2.320 0.405 ;
        RECT  0.795 1.205 2.320 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCNDD2

MACRO LNCNDD4
    CLASS CORE ;
    FOREIGN LNCNDD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.325 4.125 0.635 ;
        RECT  3.850 1.110 4.085 1.290 ;
        RECT  3.550 0.325 3.850 1.290 ;
        RECT  3.415 0.325 3.550 0.635 ;
        RECT  3.455 1.110 3.550 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.325 5.150 0.635 ;
        RECT  5.050 1.100 5.150 1.410 ;
        RECT  4.750 0.325 5.050 1.410 ;
        RECT  4.415 0.325 4.750 0.635 ;
        RECT  4.415 1.100 4.750 1.410 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.415 0.325 4.650 0.635 ;
        RECT  4.415 1.100 4.650 1.410 ;
        RECT  3.950 0.325 4.125 0.635 ;
        RECT  3.950 1.110 4.085 1.290 ;
        RECT  3.415 0.325 3.450 0.635 ;
        RECT  4.295 0.780 4.500 0.890 ;
        RECT  4.195 0.780 4.295 1.480 ;
        RECT  3.290 1.380 4.195 1.480 ;
        RECT  3.200 0.575 3.290 1.480 ;
        RECT  3.075 0.575 3.200 0.685 ;
        RECT  3.075 1.380 3.200 1.480 ;
        RECT  2.965 0.275 3.075 0.685 ;
        RECT  2.965 1.050 3.075 1.480 ;
        RECT  2.585 0.780 3.050 0.890 ;
        RECT  2.475 0.275 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.290 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.290 0.405 ;
        RECT  0.795 1.205 2.290 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.275 0.180 0.675 ;
        RECT  0.150 1.050 0.180 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LNCNDD4

MACRO LNCNDQD1
    CLASS CORE ;
    FOREIGN LNCNDQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.275 3.350 1.490 ;
        RECT  3.215 0.275 3.250 0.675 ;
        RECT  3.215 1.080 3.250 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.400 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 1.635 3.400 1.965 ;
        RECT  2.900 1.495 3.070 1.965 ;
        RECT  0.000 1.635 2.900 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.120 0.750 3.150 0.920 ;
        RECT  3.020 0.525 3.120 1.180 ;
        RECT  2.665 0.525 3.020 0.635 ;
        RECT  2.665 1.070 3.020 1.180 ;
        RECT  2.575 0.780 2.930 0.890 ;
        RECT  2.475 0.275 2.575 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.280 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.280 0.405 ;
        RECT  0.795 1.205 2.280 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCNDQD1

MACRO LNCNDQD2
    CLASS CORE ;
    FOREIGN LNCNDQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.275 3.350 1.490 ;
        RECT  3.165 0.275 3.250 0.665 ;
        RECT  3.165 1.080 3.250 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0419 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.600 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.075 0.750 3.125 0.920 ;
        RECT  2.975 0.305 3.075 1.310 ;
        RECT  2.625 0.305 2.975 0.415 ;
        RECT  2.785 1.220 2.975 1.310 ;
        RECT  2.600 0.780 2.885 0.890 ;
        RECT  2.675 1.220 2.785 1.525 ;
        RECT  2.580 0.505 2.600 0.890 ;
        RECT  2.490 0.505 2.580 1.525 ;
        RECT  2.010 1.415 2.490 1.525 ;
        RECT  2.305 0.295 2.395 1.315 ;
        RECT  1.465 0.295 2.305 0.405 ;
        RECT  0.795 1.205 2.305 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCNDQD2

MACRO LNCNDQD4
    CLASS CORE ;
    FOREIGN LNCNDQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.325 4.150 0.635 ;
        RECT  4.050 1.100 4.150 1.410 ;
        RECT  3.750 0.325 4.050 1.410 ;
        RECT  3.415 0.325 3.750 0.635 ;
        RECT  3.415 1.100 3.750 1.410 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0419 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.415 0.325 3.650 0.635 ;
        RECT  3.415 1.100 3.650 1.410 ;
        RECT  3.310 0.780 3.600 0.890 ;
        RECT  3.210 0.575 3.310 1.150 ;
        RECT  3.075 0.575 3.210 0.685 ;
        RECT  3.075 1.050 3.210 1.150 ;
        RECT  2.600 0.780 3.100 0.890 ;
        RECT  2.965 0.275 3.075 0.685 ;
        RECT  2.965 1.050 3.075 1.460 ;
        RECT  2.590 0.275 2.600 0.890 ;
        RECT  2.490 0.275 2.590 1.525 ;
        RECT  2.010 1.415 2.490 1.525 ;
        RECT  2.305 0.295 2.395 1.315 ;
        RECT  1.465 0.295 2.305 0.405 ;
        RECT  0.795 1.205 2.305 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.275 0.180 0.675 ;
        RECT  0.150 1.050 0.180 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LNCNDQD4

MACRO LNCNQD1
    CLASS CORE ;
    FOREIGN LNCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.290 3.150 1.515 ;
        RECT  2.960 0.290 3.050 0.685 ;
        RECT  2.960 1.055 3.050 1.515 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.495 ;
        RECT  1.110 1.345 1.200 1.495 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.710 0.355 1.435 ;
        RECT  0.245 0.710 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.815 -0.165 3.200 0.165 ;
        RECT  2.690 -0.165 2.815 0.465 ;
        RECT  0.000 -0.165 2.690 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.825 1.635 3.200 1.965 ;
        RECT  2.685 1.270 2.825 1.965 ;
        RECT  0.000 1.635 2.685 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.580 0.795 2.945 0.915 ;
        RECT  2.490 0.260 2.580 1.465 ;
        RECT  2.440 0.260 2.490 0.645 ;
        RECT  2.430 1.040 2.490 1.465 ;
        RECT  2.300 0.740 2.380 0.930 ;
        RECT  2.190 0.285 2.300 1.495 ;
        RECT  1.680 1.395 2.190 1.495 ;
        RECT  2.000 0.315 2.100 1.255 ;
        RECT  1.135 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.710 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.600 ;
        RECT  0.155 0.405 0.210 0.600 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.405 0.155 1.515 ;
    END
END LNCNQD1

MACRO LNCNQD2
    CLASS CORE ;
    FOREIGN LNCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.075 0.555 3.150 1.175 ;
        RECT  3.070 0.255 3.075 1.175 ;
        RECT  3.050 0.255 3.070 1.465 ;
        RECT  2.945 0.255 3.050 0.680 ;
        RECT  2.955 1.035 3.050 1.465 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.395 1.420 1.505 ;
        RECT  0.355 1.165 0.430 1.505 ;
        RECT  0.340 0.710 0.355 1.505 ;
        RECT  0.245 0.710 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.335 -0.165 3.400 0.165 ;
        RECT  3.205 -0.165 3.335 0.445 ;
        RECT  2.815 -0.165 3.205 0.165 ;
        RECT  2.700 -0.165 2.815 0.660 ;
        RECT  0.000 -0.165 2.700 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 1.635 3.400 1.965 ;
        RECT  3.210 1.310 3.330 1.965 ;
        RECT  2.815 1.635 3.210 1.965 ;
        RECT  2.700 1.045 2.815 1.965 ;
        RECT  0.000 1.635 2.700 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.610 0.770 2.940 0.900 ;
        RECT  2.510 0.305 2.610 1.485 ;
        RECT  2.395 0.305 2.510 0.405 ;
        RECT  2.440 1.270 2.510 1.485 ;
        RECT  2.330 0.740 2.420 0.930 ;
        RECT  2.230 0.495 2.330 1.505 ;
        RECT  1.680 1.395 2.230 1.505 ;
        RECT  2.005 0.315 2.110 1.255 ;
        RECT  1.130 0.315 2.005 0.405 ;
        RECT  0.540 1.165 2.005 1.255 ;
        RECT  1.340 0.985 1.710 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.600 ;
        RECT  0.155 0.405 0.210 0.600 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.405 0.155 1.515 ;
    END
END LNCNQD2

MACRO LNCNQD4
    CLASS CORE ;
    FOREIGN LNCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 0.310 3.860 0.690 ;
        RECT  3.750 1.110 3.860 1.490 ;
        RECT  3.650 0.545 3.750 0.690 ;
        RECT  3.650 1.110 3.750 1.210 ;
        RECT  3.350 0.545 3.650 1.210 ;
        RECT  3.240 0.310 3.350 0.690 ;
        RECT  3.345 1.110 3.350 1.210 ;
        RECT  3.240 1.110 3.345 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0812 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.425 1.415 1.400 1.525 ;
        RECT  0.355 1.175 0.425 1.525 ;
        RECT  0.335 0.700 0.355 1.525 ;
        RECT  0.240 0.700 0.335 1.265 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0406 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.495 1.875 0.665 ;
        RECT  1.445 0.495 1.555 0.890 ;
        RECT  0.750 0.495 1.445 0.585 ;
        RECT  0.650 0.255 0.750 0.585 ;
        RECT  0.440 0.255 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.690 ;
        RECT  3.605 -0.165 4.015 0.165 ;
        RECT  3.495 -0.165 3.605 0.455 ;
        RECT  3.085 -0.165 3.495 0.165 ;
        RECT  2.975 -0.165 3.085 0.690 ;
        RECT  2.605 -0.165 2.975 0.165 ;
        RECT  2.415 -0.165 2.605 0.445 ;
        RECT  0.000 -0.165 2.415 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.110 4.125 1.965 ;
        RECT  3.605 1.635 4.015 1.965 ;
        RECT  3.495 1.320 3.605 1.965 ;
        RECT  3.085 1.635 3.495 1.965 ;
        RECT  2.975 1.110 3.085 1.965 ;
        RECT  2.565 1.635 2.975 1.965 ;
        RECT  2.455 1.320 2.565 1.965 ;
        RECT  0.000 1.635 2.455 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 0.310 3.860 0.690 ;
        RECT  3.750 1.110 3.860 1.490 ;
        RECT  3.240 0.310 3.250 0.690 ;
        RECT  3.240 1.110 3.250 1.490 ;
        RECT  2.825 0.800 3.260 0.910 ;
        RECT  2.715 0.310 2.825 1.490 ;
        RECT  2.400 0.555 2.510 1.230 ;
        RECT  2.255 0.555 2.400 0.690 ;
        RECT  2.255 1.110 2.400 1.230 ;
        RECT  2.145 0.310 2.255 0.690 ;
        RECT  2.145 1.110 2.255 1.525 ;
        RECT  1.660 1.415 2.145 1.525 ;
        RECT  2.055 0.775 2.100 0.945 ;
        RECT  1.965 0.315 2.055 1.305 ;
        RECT  1.115 0.315 1.965 0.405 ;
        RECT  0.515 1.195 1.965 1.305 ;
        RECT  1.355 1.000 1.690 1.105 ;
        RECT  1.245 0.675 1.355 1.105 ;
        RECT  1.040 0.675 1.245 0.785 ;
        RECT  0.555 0.985 1.245 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.205 0.495 0.445 0.585 ;
        RECT  0.150 1.355 0.225 1.525 ;
        RECT  0.150 0.390 0.205 0.585 ;
        RECT  0.060 0.390 0.150 1.525 ;
    END
END LNCNQD4

MACRO LNCSND1
    CLASS CORE ;
    FOREIGN LNCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.710 2.370 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.155 3.290 1.255 ;
        RECT  3.150 0.295 3.255 0.670 ;
        RECT  3.135 0.295 3.150 1.255 ;
        RECT  3.050 0.510 3.135 1.255 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 0.285 3.750 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.495 ;
        RECT  1.110 1.345 1.200 1.495 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.710 0.355 1.435 ;
        RECT  0.245 0.710 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.380 0.730 3.490 1.500 ;
        RECT  2.915 1.380 3.380 1.500 ;
        RECT  2.815 0.305 2.915 1.500 ;
        RECT  2.590 0.305 2.815 0.420 ;
        RECT  2.590 1.380 2.815 1.500 ;
        RECT  2.595 0.510 2.705 1.270 ;
        RECT  2.330 0.510 2.595 0.600 ;
        RECT  2.480 1.180 2.595 1.270 ;
        RECT  2.390 1.180 2.480 1.495 ;
        RECT  1.680 1.395 2.390 1.495 ;
        RECT  2.000 0.315 2.115 1.255 ;
        RECT  1.130 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.700 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.600 ;
        RECT  0.155 0.405 0.210 0.600 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.405 0.155 1.515 ;
    END
END LNCSND1

MACRO LNCSND2
    CLASS CORE ;
    FOREIGN LNCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.510 2.370 0.940 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.230 0.275 3.350 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.865 0.510 3.950 1.195 ;
        RECT  3.850 0.275 3.865 1.490 ;
        RECT  3.755 0.275 3.850 0.675 ;
        RECT  3.755 1.045 3.850 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.495 ;
        RECT  1.110 1.345 1.200 1.495 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.710 0.355 1.435 ;
        RECT  0.245 0.710 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.445 ;
        RECT  3.615 -0.165 4.015 0.165 ;
        RECT  3.490 -0.165 3.615 0.675 ;
        RECT  3.095 -0.165 3.490 0.165 ;
        RECT  2.970 -0.165 3.095 0.675 ;
        RECT  0.000 -0.165 2.970 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 1.635 4.200 1.965 ;
        RECT  4.010 1.325 4.130 1.965 ;
        RECT  2.540 1.635 4.010 1.965 ;
        RECT  2.435 1.310 2.540 1.965 ;
        RECT  0.000 1.635 2.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.785 3.760 0.885 ;
        RECT  3.495 0.785 3.605 1.505 ;
        RECT  2.830 1.395 3.495 1.505 ;
        RECT  2.710 0.270 2.830 1.505 ;
        RECT  2.510 0.330 2.620 1.190 ;
        RECT  2.330 0.330 2.510 0.420 ;
        RECT  2.325 1.100 2.510 1.190 ;
        RECT  2.235 1.100 2.325 1.495 ;
        RECT  1.680 1.395 2.235 1.495 ;
        RECT  2.000 0.315 2.115 1.255 ;
        RECT  1.135 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.710 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.600 ;
        RECT  0.155 0.405 0.210 0.600 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.405 0.155 1.515 ;
    END
END LNCSND2

MACRO LNCSND4
    CLASS CORE ;
    FOREIGN LNCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.700 2.550 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.310 4.305 0.695 ;
        RECT  4.050 1.110 4.305 1.290 ;
        RECT  3.750 0.310 4.050 1.290 ;
        RECT  3.615 0.310 3.750 0.695 ;
        RECT  3.615 1.110 3.750 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.310 5.305 0.690 ;
        RECT  5.250 1.110 5.305 1.490 ;
        RECT  4.950 0.310 5.250 1.490 ;
        RECT  4.615 0.310 4.950 0.690 ;
        RECT  4.615 1.110 4.950 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.505 ;
        RECT  1.110 1.345 1.200 1.505 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.700 0.355 1.435 ;
        RECT  0.245 0.700 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.525 -0.165 5.600 0.165 ;
        RECT  5.415 -0.165 5.525 0.690 ;
        RECT  0.000 -0.165 5.415 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.525 1.635 5.600 1.965 ;
        RECT  5.415 1.110 5.525 1.965 ;
        RECT  0.000 1.635 5.415 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.615 0.310 4.850 0.690 ;
        RECT  4.615 1.110 4.850 1.490 ;
        RECT  4.150 0.310 4.305 0.695 ;
        RECT  4.150 1.110 4.305 1.290 ;
        RECT  3.615 0.310 3.650 0.695 ;
        RECT  3.615 1.110 3.650 1.290 ;
        RECT  4.505 0.800 4.750 0.910 ;
        RECT  4.415 0.800 4.505 1.505 ;
        RECT  3.265 1.400 4.415 1.505 ;
        RECT  3.370 0.600 3.480 1.200 ;
        RECT  3.265 0.600 3.370 0.690 ;
        RECT  3.265 1.110 3.370 1.200 ;
        RECT  3.155 0.310 3.265 0.690 ;
        RECT  3.155 1.110 3.265 1.505 ;
        RECT  3.065 0.800 3.260 0.910 ;
        RECT  2.955 0.345 3.065 1.505 ;
        RECT  2.355 0.345 2.955 0.455 ;
        RECT  1.680 1.395 2.955 1.505 ;
        RECT  2.735 0.700 2.845 1.285 ;
        RECT  2.115 1.180 2.735 1.285 ;
        RECT  2.000 0.315 2.115 1.285 ;
        RECT  1.135 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.710 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.585 ;
        RECT  0.155 0.390 0.210 0.585 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.390 0.155 1.515 ;
    END
END LNCSND4

MACRO LNCSNDD1
    CLASS CORE ;
    FOREIGN LNCSNDD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.750 1.090 ;
        RECT  2.630 0.710 2.650 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 1.015 3.655 1.125 ;
        RECT  3.550 0.275 3.605 0.675 ;
        RECT  3.450 0.275 3.550 1.125 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.275 4.150 1.490 ;
        RECT  4.025 0.275 4.050 0.675 ;
        RECT  4.015 1.080 4.050 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.865 -0.165 4.200 0.165 ;
        RECT  3.755 -0.165 3.865 0.655 ;
        RECT  3.070 -0.165 3.755 0.165 ;
        RECT  2.960 -0.165 3.070 0.355 ;
        RECT  0.880 -0.165 2.960 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.895 1.635 4.200 1.965 ;
        RECT  3.725 1.395 3.895 1.965 ;
        RECT  3.030 1.635 3.725 1.965 ;
        RECT  2.860 1.495 3.030 1.965 ;
        RECT  0.000 1.635 2.860 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.870 0.750 3.950 0.920 ;
        RECT  3.770 0.750 3.870 1.305 ;
        RECT  3.355 1.215 3.770 1.305 ;
        RECT  3.245 0.275 3.355 1.460 ;
        RECT  3.025 0.490 3.135 1.300 ;
        RECT  2.675 0.490 3.025 0.600 ;
        RECT  2.645 1.200 3.025 1.300 ;
        RECT  2.535 1.200 2.645 1.525 ;
        RECT  2.010 1.415 2.535 1.525 ;
        RECT  2.380 0.750 2.480 0.920 ;
        RECT  2.280 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.280 0.405 ;
        RECT  0.795 1.205 2.280 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCSNDD1

MACRO LNCSNDD2
    CLASS CORE ;
    FOREIGN LNCSNDD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.750 2.670 0.920 ;
        RECT  2.550 0.600 2.615 0.920 ;
        RECT  2.525 0.310 2.550 0.920 ;
        RECT  2.450 0.310 2.525 0.690 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.275 3.565 1.180 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.065 0.585 4.150 1.150 ;
        RECT  4.050 0.275 4.065 1.460 ;
        RECT  3.955 0.275 4.050 0.685 ;
        RECT  3.955 1.050 4.050 1.460 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.485 ;
        RECT  0.880 -0.165 4.215 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.250 4.325 1.965 ;
        RECT  0.000 1.635 4.215 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.820 0.780 3.960 0.890 ;
        RECT  3.720 0.780 3.820 1.370 ;
        RECT  3.295 1.270 3.720 1.370 ;
        RECT  3.195 0.575 3.295 1.370 ;
        RECT  3.065 0.575 3.195 0.685 ;
        RECT  3.065 1.270 3.195 1.370 ;
        RECT  2.865 0.780 3.095 0.890 ;
        RECT  2.955 0.275 3.065 0.685 ;
        RECT  2.955 1.050 3.065 1.460 ;
        RECT  2.815 0.575 2.865 1.150 ;
        RECT  2.775 0.275 2.815 1.150 ;
        RECT  2.705 0.275 2.775 0.665 ;
        RECT  2.585 1.050 2.775 1.150 ;
        RECT  2.475 1.050 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.350 0.780 2.430 0.890 ;
        RECT  2.260 0.295 2.350 1.315 ;
        RECT  1.465 0.295 2.260 0.405 ;
        RECT  0.795 1.205 2.260 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCSNDD2

MACRO LNCSNDD4
    CLASS CORE ;
    FOREIGN LNCSNDD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.700 2.760 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.325 4.665 0.635 ;
        RECT  4.450 1.110 4.655 1.290 ;
        RECT  4.150 0.325 4.450 1.290 ;
        RECT  3.945 0.325 4.150 0.635 ;
        RECT  3.955 1.110 4.150 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.325 5.685 0.635 ;
        RECT  5.650 1.100 5.685 1.410 ;
        RECT  5.350 0.325 5.650 1.410 ;
        RECT  4.965 0.325 5.350 0.635 ;
        RECT  4.965 1.100 5.350 1.410 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.895 -0.165 6.000 0.165 ;
        RECT  5.785 -0.165 5.895 0.685 ;
        RECT  0.000 -0.165 5.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.895 1.635 6.000 1.965 ;
        RECT  5.785 1.050 5.895 1.965 ;
        RECT  0.000 1.635 5.785 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.965 0.325 5.250 0.635 ;
        RECT  4.965 1.100 5.250 1.410 ;
        RECT  4.550 0.325 4.665 0.635 ;
        RECT  4.550 1.110 4.655 1.290 ;
        RECT  3.945 0.325 4.050 0.635 ;
        RECT  3.955 1.110 4.050 1.290 ;
        RECT  4.865 0.780 5.110 0.890 ;
        RECT  4.775 0.780 4.865 1.505 ;
        RECT  3.595 1.400 4.775 1.505 ;
        RECT  3.735 0.600 3.835 1.195 ;
        RECT  3.595 0.600 3.735 0.690 ;
        RECT  3.595 1.095 3.735 1.195 ;
        RECT  3.485 0.310 3.595 0.690 ;
        RECT  3.485 1.095 3.595 1.505 ;
        RECT  3.395 0.780 3.590 0.890 ;
        RECT  3.295 0.490 3.395 1.495 ;
        RECT  2.675 0.490 3.295 0.600 ;
        RECT  2.525 1.385 3.295 1.495 ;
        RECT  3.070 0.750 3.180 1.285 ;
        RECT  2.420 1.180 3.070 1.285 ;
        RECT  2.415 1.385 2.525 1.525 ;
        RECT  2.310 0.295 2.420 1.285 ;
        RECT  2.010 1.415 2.415 1.525 ;
        RECT  1.465 0.295 2.310 0.405 ;
        RECT  2.230 1.180 2.310 1.285 ;
        RECT  2.130 1.180 2.230 1.315 ;
        RECT  0.795 1.205 2.130 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.275 0.180 0.675 ;
        RECT  0.150 1.050 0.180 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LNCSNDD4

MACRO LNCSNDQD1
    CLASS CORE ;
    FOREIGN LNCSNDQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.770 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.275 3.550 1.490 ;
        RECT  3.415 0.275 3.450 0.675 ;
        RECT  3.415 1.080 3.450 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.600 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.305 0.750 3.360 0.920 ;
        RECT  3.205 0.310 3.305 1.145 ;
        RECT  2.865 0.310 3.205 0.420 ;
        RECT  2.865 1.035 3.205 1.145 ;
        RECT  2.985 0.510 3.095 0.930 ;
        RECT  2.560 0.510 2.985 0.620 ;
        RECT  2.560 1.250 2.575 1.525 ;
        RECT  2.470 0.510 2.560 1.525 ;
        RECT  2.010 1.415 2.470 1.525 ;
        RECT  2.280 0.295 2.380 1.315 ;
        RECT  1.465 0.295 2.280 0.405 ;
        RECT  0.795 1.205 2.280 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCSNDQD1

MACRO LNCSNDQD2
    CLASS CORE ;
    FOREIGN LNCSNDQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.750 2.670 0.920 ;
        RECT  2.550 0.600 2.615 0.920 ;
        RECT  2.525 0.310 2.550 0.920 ;
        RECT  2.450 0.310 2.525 0.690 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.585 3.750 1.150 ;
        RECT  3.615 0.585 3.650 0.685 ;
        RECT  3.615 1.050 3.650 1.150 ;
        RECT  3.505 0.275 3.615 0.685 ;
        RECT  3.505 1.050 3.615 1.460 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.875 -0.165 4.000 0.165 ;
        RECT  3.765 -0.165 3.875 0.475 ;
        RECT  3.365 -0.165 3.765 0.165 ;
        RECT  3.245 -0.165 3.365 0.475 ;
        RECT  0.880 -0.165 3.245 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.875 1.635 4.000 1.965 ;
        RECT  3.765 1.250 3.875 1.965 ;
        RECT  3.365 1.635 3.765 1.965 ;
        RECT  3.245 1.250 3.365 1.965 ;
        RECT  2.845 1.635 3.245 1.965 ;
        RECT  2.735 1.250 2.845 1.965 ;
        RECT  0.000 1.635 2.735 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.325 0.780 3.540 0.890 ;
        RECT  3.225 0.575 3.325 1.150 ;
        RECT  3.095 0.575 3.225 0.685 ;
        RECT  3.095 1.050 3.225 1.150 ;
        RECT  2.865 0.780 3.125 0.890 ;
        RECT  2.985 0.275 3.095 0.685 ;
        RECT  2.985 1.050 3.095 1.460 ;
        RECT  2.815 0.575 2.865 1.150 ;
        RECT  2.775 0.275 2.815 1.150 ;
        RECT  2.705 0.275 2.775 0.665 ;
        RECT  2.585 1.050 2.775 1.150 ;
        RECT  2.475 1.050 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.350 0.780 2.430 0.890 ;
        RECT  2.260 0.295 2.350 1.315 ;
        RECT  1.465 0.295 2.260 0.405 ;
        RECT  0.795 1.205 2.260 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNCSNDQD2

MACRO LNCSNDQD4
    CLASS CORE ;
    FOREIGN LNCSNDQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.750 1.090 ;
        RECT  2.570 0.710 2.650 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.325 4.350 0.635 ;
        RECT  4.250 1.100 4.350 1.410 ;
        RECT  3.950 0.325 4.250 1.410 ;
        RECT  3.615 0.325 3.950 0.635 ;
        RECT  3.615 1.100 3.950 1.410 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0474 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0420 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.495 2.170 0.690 ;
        RECT  0.950 0.495 2.060 0.585 ;
        RECT  0.840 0.495 0.950 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.960 1.635 4.600 1.965 ;
        RECT  2.790 1.390 2.960 1.965 ;
        RECT  0.000 1.635 2.790 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.615 0.325 3.850 0.635 ;
        RECT  3.615 1.100 3.850 1.410 ;
        RECT  3.505 0.780 3.770 0.890 ;
        RECT  3.405 0.575 3.505 1.150 ;
        RECT  3.275 0.575 3.405 0.685 ;
        RECT  3.275 1.050 3.405 1.150 ;
        RECT  2.960 0.780 3.305 0.890 ;
        RECT  3.165 0.275 3.275 0.685 ;
        RECT  3.165 1.050 3.275 1.460 ;
        RECT  2.860 0.490 2.960 1.300 ;
        RECT  2.635 0.490 2.860 0.600 ;
        RECT  2.585 1.200 2.860 1.300 ;
        RECT  2.475 1.200 2.585 1.525 ;
        RECT  2.010 1.415 2.475 1.525 ;
        RECT  2.350 0.750 2.420 0.920 ;
        RECT  2.260 0.295 2.350 1.315 ;
        RECT  1.465 0.295 2.260 0.405 ;
        RECT  0.795 1.205 2.260 1.315 ;
        RECT  1.550 0.995 2.020 1.105 ;
        RECT  1.535 1.435 1.745 1.545 ;
        RECT  1.440 0.675 1.550 1.105 ;
        RECT  0.180 1.435 1.535 1.525 ;
        RECT  0.685 1.015 1.440 1.105 ;
        RECT  0.360 0.490 0.715 0.600 ;
        RECT  0.575 1.015 0.685 1.340 ;
        RECT  0.360 1.015 0.575 1.105 ;
        RECT  0.270 0.490 0.360 1.105 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.275 0.180 0.675 ;
        RECT  0.150 1.050 0.180 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LNCSNDQD4

MACRO LNCSNQD1
    CLASS CORE ;
    FOREIGN LNCSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.510 2.370 1.065 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.275 3.350 1.515 ;
        RECT  3.215 0.275 3.250 0.680 ;
        RECT  3.215 1.030 3.250 1.515 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.495 ;
        RECT  1.110 1.345 1.200 1.495 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.710 0.355 1.435 ;
        RECT  0.245 0.710 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.165 3.400 0.165 ;
        RECT  2.945 -0.165 3.070 0.465 ;
        RECT  0.000 -0.165 2.945 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.635 3.400 1.965 ;
        RECT  2.940 1.270 3.080 1.965 ;
        RECT  2.535 1.635 2.940 1.965 ;
        RECT  2.425 1.355 2.535 1.965 ;
        RECT  0.000 1.635 2.425 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.820 0.765 3.140 0.935 ;
        RECT  2.720 0.260 2.820 1.480 ;
        RECT  2.695 0.260 2.720 0.645 ;
        RECT  2.695 1.040 2.720 1.480 ;
        RECT  2.595 0.750 2.620 0.920 ;
        RECT  2.480 0.330 2.595 1.265 ;
        RECT  2.330 0.330 2.480 0.420 ;
        RECT  2.310 1.175 2.480 1.265 ;
        RECT  2.220 1.175 2.310 1.495 ;
        RECT  1.680 1.395 2.220 1.495 ;
        RECT  2.000 0.315 2.115 1.255 ;
        RECT  1.145 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.710 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.600 ;
        RECT  0.155 0.405 0.210 0.600 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.405 0.155 1.515 ;
    END
END LNCSNQD1

MACRO LNCSNQD2
    CLASS CORE ;
    FOREIGN LNCSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.650 2.370 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.275 0.540 3.350 1.195 ;
        RECT  3.250 0.275 3.275 1.490 ;
        RECT  3.145 0.275 3.250 0.655 ;
        RECT  3.145 1.045 3.250 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0538 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.495 ;
        RECT  1.110 1.345 1.200 1.495 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.710 0.355 1.435 ;
        RECT  0.245 0.710 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 -0.165 3.600 0.165 ;
        RECT  3.405 -0.165 3.535 0.445 ;
        RECT  0.000 -0.165 3.405 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 1.635 3.600 1.965 ;
        RECT  3.405 1.315 3.535 1.965 ;
        RECT  0.000 1.635 3.405 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.830 0.750 3.130 0.920 ;
        RECT  2.730 0.270 2.830 1.505 ;
        RECT  2.645 0.270 2.730 0.655 ;
        RECT  2.645 1.045 2.730 1.505 ;
        RECT  2.555 0.750 2.620 0.940 ;
        RECT  2.465 0.330 2.555 1.495 ;
        RECT  2.330 0.330 2.465 0.420 ;
        RECT  1.680 1.395 2.465 1.495 ;
        RECT  2.000 0.315 2.115 1.255 ;
        RECT  1.135 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.700 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.600 ;
        RECT  0.155 0.405 0.210 0.600 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.405 0.155 1.515 ;
    END
END LNCSNQD2

MACRO LNCSNQD4
    CLASS CORE ;
    FOREIGN LNCSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.510 2.370 0.940 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.740 0.295 3.875 0.690 ;
        RECT  3.745 1.020 3.875 1.515 ;
        RECT  3.670 1.020 3.745 1.200 ;
        RECT  3.670 0.510 3.740 0.690 ;
        RECT  3.355 0.510 3.670 1.200 ;
        RECT  3.350 0.295 3.355 1.515 ;
        RECT  3.225 0.295 3.350 0.690 ;
        RECT  3.225 1.020 3.350 1.515 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.395 1.420 1.495 ;
        RECT  1.110 1.345 1.200 1.495 ;
        RECT  0.430 1.345 1.110 1.435 ;
        RECT  0.355 1.165 0.430 1.435 ;
        RECT  0.340 0.700 0.355 1.435 ;
        RECT  0.245 0.700 0.340 1.255 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0380 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0405 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.890 0.645 ;
        RECT  1.450 0.495 1.550 0.890 ;
        RECT  0.750 0.495 1.450 0.585 ;
        RECT  0.650 0.275 0.750 0.585 ;
        RECT  0.480 0.275 0.650 0.385 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.005 -0.165 4.125 0.690 ;
        RECT  3.635 -0.165 4.005 0.165 ;
        RECT  3.465 -0.165 3.635 0.420 ;
        RECT  3.095 -0.165 3.465 0.165 ;
        RECT  2.965 -0.165 3.095 0.675 ;
        RECT  0.000 -0.165 2.965 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.135 1.635 4.200 1.965 ;
        RECT  4.015 1.095 4.135 1.965 ;
        RECT  3.615 1.635 4.015 1.965 ;
        RECT  3.485 1.310 3.615 1.965 ;
        RECT  3.085 1.635 3.485 1.965 ;
        RECT  2.975 1.060 3.085 1.965 ;
        RECT  2.565 1.635 2.975 1.965 ;
        RECT  2.425 1.310 2.565 1.965 ;
        RECT  0.000 1.635 2.425 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 0.295 3.875 0.690 ;
        RECT  3.750 1.020 3.875 1.515 ;
        RECT  3.225 0.295 3.250 0.690 ;
        RECT  3.225 1.020 3.250 1.515 ;
        RECT  2.830 0.790 3.220 0.900 ;
        RECT  2.720 0.270 2.830 1.525 ;
        RECT  2.490 0.330 2.620 1.190 ;
        RECT  2.330 0.330 2.490 0.420 ;
        RECT  2.325 1.100 2.490 1.190 ;
        RECT  2.225 1.100 2.325 1.495 ;
        RECT  1.680 1.395 2.225 1.495 ;
        RECT  2.000 0.315 2.115 1.255 ;
        RECT  1.135 0.315 2.000 0.405 ;
        RECT  0.540 1.165 2.000 1.255 ;
        RECT  1.340 0.985 1.710 1.075 ;
        RECT  1.250 0.675 1.340 1.075 ;
        RECT  1.060 0.675 1.250 0.765 ;
        RECT  0.555 0.985 1.250 1.075 ;
        RECT  0.445 0.495 0.555 1.075 ;
        RECT  0.210 0.495 0.445 0.585 ;
        RECT  0.155 0.390 0.210 0.585 ;
        RECT  0.155 1.345 0.210 1.515 ;
        RECT  0.065 0.390 0.155 1.515 ;
    END
END LNCSNQD4

MACRO LND1
    CLASS CORE ;
    FOREIGN LND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.275 2.950 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.545 2.555 1.290 ;
        RECT  2.400 0.545 2.445 0.675 ;
        RECT  2.290 1.110 2.445 1.290 ;
        RECT  2.290 0.275 2.400 0.675 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.095 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.895 -0.165 3.000 0.165 ;
        RECT  1.745 -0.165 1.895 0.455 ;
        RECT  0.000 -0.165 1.745 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.635 3.000 1.965 ;
        RECT  0.950 1.205 1.040 1.965 ;
        RECT  0.805 1.205 0.950 1.305 ;
        RECT  0.000 1.635 0.950 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.645 0.730 2.735 1.490 ;
        RECT  2.200 1.400 2.645 1.490 ;
        RECT  2.110 0.275 2.200 1.490 ;
        RECT  2.030 0.275 2.110 0.645 ;
        RECT  2.030 1.245 2.110 1.490 ;
        RECT  1.770 0.545 2.030 0.645 ;
        RECT  1.910 0.755 2.020 1.135 ;
        RECT  1.540 1.045 1.910 1.135 ;
        RECT  1.660 0.545 1.770 0.935 ;
        RECT  1.220 1.435 1.550 1.525 ;
        RECT  1.440 0.275 1.540 1.135 ;
        RECT  1.310 0.275 1.440 0.475 ;
        RECT  1.420 1.045 1.440 1.135 ;
        RECT  1.310 1.045 1.420 1.345 ;
        RECT  1.220 0.575 1.350 0.685 ;
        RECT  1.130 0.305 1.220 1.525 ;
        RECT  0.410 0.305 1.130 0.405 ;
        RECT  0.715 1.415 0.860 1.525 ;
        RECT  0.610 0.495 0.715 1.525 ;
        RECT  0.535 0.495 0.610 0.615 ;
        RECT  0.580 1.060 0.610 1.525 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.305 0.410 1.310 ;
        RECT  0.065 0.305 0.310 0.495 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LND1

MACRO LND2
    CLASS CORE ;
    FOREIGN LND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.150 1.490 ;
        RECT  2.965 0.275 3.050 0.675 ;
        RECT  2.965 1.055 3.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.275 2.595 1.290 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.095 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.635 3.400 1.965 ;
        RECT  0.950 1.205 1.040 1.965 ;
        RECT  0.805 1.205 0.950 1.305 ;
        RECT  0.000 1.635 0.950 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.855 0.790 2.955 0.890 ;
        RECT  2.755 0.790 2.855 1.490 ;
        RECT  2.175 1.400 2.755 1.490 ;
        RECT  2.085 0.275 2.175 1.490 ;
        RECT  1.995 0.275 2.085 0.645 ;
        RECT  1.995 1.245 2.085 1.490 ;
        RECT  1.755 0.545 1.995 0.645 ;
        RECT  1.885 0.755 1.995 1.135 ;
        RECT  1.520 1.045 1.885 1.135 ;
        RECT  1.645 0.545 1.755 0.935 ;
        RECT  1.220 1.435 1.545 1.525 ;
        RECT  1.420 0.275 1.520 1.135 ;
        RECT  1.310 0.275 1.420 0.475 ;
        RECT  1.310 1.045 1.420 1.345 ;
        RECT  1.220 0.575 1.330 0.685 ;
        RECT  1.130 0.305 1.220 1.525 ;
        RECT  0.410 0.305 1.130 0.405 ;
        RECT  0.715 1.415 0.860 1.525 ;
        RECT  0.610 0.495 0.715 1.525 ;
        RECT  0.535 0.495 0.610 0.615 ;
        RECT  0.580 1.060 0.610 1.525 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.305 0.410 1.310 ;
        RECT  0.065 0.305 0.310 0.495 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LND2

MACRO LND4
    CLASS CORE ;
    FOREIGN LND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.310 4.150 0.690 ;
        RECT  4.050 1.110 4.150 1.490 ;
        RECT  3.750 0.310 4.050 1.490 ;
        RECT  3.425 0.310 3.750 0.690 ;
        RECT  3.425 1.110 3.750 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.150 0.690 ;
        RECT  3.050 1.110 3.115 1.290 ;
        RECT  2.750 0.310 3.050 1.290 ;
        RECT  2.425 0.310 2.750 0.690 ;
        RECT  2.425 1.110 2.750 1.290 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.095 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.635 4.400 1.965 ;
        RECT  0.950 1.205 1.040 1.965 ;
        RECT  0.805 1.205 0.950 1.305 ;
        RECT  0.000 1.635 0.950 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.425 0.310 3.650 0.690 ;
        RECT  3.425 1.110 3.650 1.490 ;
        RECT  2.425 0.310 2.650 0.690 ;
        RECT  2.425 1.110 2.650 1.290 ;
        RECT  3.335 0.790 3.550 0.890 ;
        RECT  3.235 0.790 3.335 1.490 ;
        RECT  2.175 1.400 3.235 1.490 ;
        RECT  2.085 0.275 2.175 1.490 ;
        RECT  1.995 0.275 2.085 0.645 ;
        RECT  1.995 1.245 2.085 1.490 ;
        RECT  1.755 0.545 1.995 0.645 ;
        RECT  1.885 0.755 1.995 1.135 ;
        RECT  1.520 1.045 1.885 1.135 ;
        RECT  1.645 0.545 1.755 0.935 ;
        RECT  1.220 1.435 1.545 1.525 ;
        RECT  1.420 0.275 1.520 1.135 ;
        RECT  1.310 0.275 1.420 0.475 ;
        RECT  1.310 1.045 1.420 1.345 ;
        RECT  1.220 0.575 1.330 0.685 ;
        RECT  1.130 0.305 1.220 1.525 ;
        RECT  0.410 0.305 1.130 0.405 ;
        RECT  0.715 1.415 0.860 1.525 ;
        RECT  0.610 0.495 0.715 1.525 ;
        RECT  0.535 0.495 0.610 0.615 ;
        RECT  0.580 1.060 0.610 1.525 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.305 0.410 1.310 ;
        RECT  0.065 0.305 0.310 0.495 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LND4

MACRO LNQD1
    CLASS CORE ;
    FOREIGN LNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.275 2.750 1.505 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.095 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.165 2.800 0.165 ;
        RECT  2.315 -0.165 2.430 0.705 ;
        RECT  1.895 -0.165 2.315 0.165 ;
        RECT  1.765 -0.165 1.895 0.455 ;
        RECT  0.000 -0.165 1.765 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.635 2.800 1.965 ;
        RECT  2.315 1.035 2.430 1.965 ;
        RECT  1.900 1.635 2.315 1.965 ;
        RECT  1.790 1.155 1.900 1.965 ;
        RECT  1.040 1.635 1.790 1.965 ;
        RECT  0.950 1.205 1.040 1.965 ;
        RECT  0.805 1.205 0.950 1.305 ;
        RECT  0.000 1.635 0.950 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.135 0.275 2.225 1.305 ;
        RECT  2.055 0.275 2.135 0.645 ;
        RECT  2.010 1.195 2.135 1.305 ;
        RECT  1.770 0.545 2.055 0.645 ;
        RECT  1.935 0.755 2.045 1.065 ;
        RECT  1.540 0.975 1.935 1.065 ;
        RECT  1.660 0.545 1.770 0.885 ;
        RECT  1.440 0.275 1.540 1.065 ;
        RECT  1.220 1.435 1.540 1.525 ;
        RECT  1.310 0.975 1.420 1.345 ;
        RECT  1.220 0.575 1.350 0.685 ;
        RECT  1.130 0.305 1.220 1.525 ;
        RECT  0.410 0.305 1.130 0.405 ;
        RECT  0.715 1.415 0.860 1.525 ;
        RECT  0.610 0.495 0.715 1.525 ;
        RECT  0.535 0.495 0.610 0.615 ;
        RECT  0.580 1.060 0.610 1.525 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.305 0.410 1.310 ;
        RECT  0.065 0.305 0.310 0.495 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
        RECT  1.310 0.275 1.440 0.475 ;
        RECT  1.420 0.975 1.440 1.065 ;
    END
END LNQD1

MACRO LNQD2
    CLASS CORE ;
    FOREIGN LNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.675 0.565 2.755 1.145 ;
        RECT  2.645 0.265 2.675 1.515 ;
        RECT  2.545 0.265 2.645 0.695 ;
        RECT  2.545 1.035 2.645 1.515 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0287 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.095 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.935 -0.165 3.000 0.165 ;
        RECT  2.805 -0.165 2.935 0.465 ;
        RECT  2.415 -0.165 2.805 0.165 ;
        RECT  2.295 -0.165 2.415 0.705 ;
        RECT  1.905 -0.165 2.295 0.165 ;
        RECT  1.750 -0.165 1.905 0.445 ;
        RECT  0.000 -0.165 1.750 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.935 1.635 3.000 1.965 ;
        RECT  2.805 1.300 2.935 1.965 ;
        RECT  2.415 1.635 2.805 1.965 ;
        RECT  2.295 1.035 2.415 1.965 ;
        RECT  1.885 1.635 2.295 1.965 ;
        RECT  1.775 1.155 1.885 1.965 ;
        RECT  1.040 1.635 1.775 1.965 ;
        RECT  0.950 1.205 1.040 1.965 ;
        RECT  0.805 1.205 0.950 1.305 ;
        RECT  0.000 1.635 0.950 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.105 0.275 2.205 1.305 ;
        RECT  2.040 0.275 2.105 0.645 ;
        RECT  1.995 1.195 2.105 1.305 ;
        RECT  1.755 0.545 2.040 0.645 ;
        RECT  1.905 0.755 2.015 1.065 ;
        RECT  1.520 0.975 1.905 1.065 ;
        RECT  1.645 0.545 1.755 0.885 ;
        RECT  1.220 1.435 1.545 1.525 ;
        RECT  1.420 0.275 1.520 1.065 ;
        RECT  1.310 0.275 1.420 0.475 ;
        RECT  1.310 0.975 1.420 1.345 ;
        RECT  1.220 0.575 1.330 0.685 ;
        RECT  1.130 0.305 1.220 1.525 ;
        RECT  0.410 0.305 1.130 0.405 ;
        RECT  0.715 1.415 0.860 1.525 ;
        RECT  0.610 0.495 0.715 1.525 ;
        RECT  0.535 0.495 0.610 0.615 ;
        RECT  0.580 1.060 0.610 1.525 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.305 0.410 1.310 ;
        RECT  0.065 0.305 0.310 0.495 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LNQD2

MACRO LNQD4
    CLASS CORE ;
    FOREIGN LNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.830 0.345 3.125 0.635 ;
        RECT  2.830 1.095 3.125 1.385 ;
        RECT  2.550 0.345 2.830 1.385 ;
        RECT  2.415 0.345 2.550 0.635 ;
        RECT  2.415 1.095 2.550 1.385 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.700 0.955 1.095 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.635 3.400 1.965 ;
        RECT  0.950 1.205 1.040 1.965 ;
        RECT  0.805 1.205 0.950 1.305 ;
        RECT  0.000 1.635 0.950 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.345 3.125 0.635 ;
        RECT  2.950 1.095 3.125 1.385 ;
        RECT  2.415 0.345 2.450 0.635 ;
        RECT  2.415 1.095 2.450 1.385 ;
        RECT  2.115 0.545 2.225 1.370 ;
        RECT  1.980 0.275 2.115 0.645 ;
        RECT  2.105 1.245 2.115 1.370 ;
        RECT  1.980 1.245 2.105 1.490 ;
        RECT  1.895 0.755 2.005 1.135 ;
        RECT  1.755 0.545 1.980 0.645 ;
        RECT  1.520 1.045 1.895 1.135 ;
        RECT  1.645 0.545 1.755 0.935 ;
        RECT  1.220 1.435 1.545 1.525 ;
        RECT  1.420 0.275 1.520 1.135 ;
        RECT  1.310 0.275 1.420 0.475 ;
        RECT  1.310 1.045 1.420 1.345 ;
        RECT  1.220 0.575 1.330 0.685 ;
        RECT  1.130 0.305 1.220 1.525 ;
        RECT  0.410 0.305 1.130 0.405 ;
        RECT  0.715 1.415 0.860 1.525 ;
        RECT  0.610 0.495 0.715 1.525 ;
        RECT  0.535 0.495 0.610 0.615 ;
        RECT  0.580 1.060 0.610 1.525 ;
        RECT  0.410 0.725 0.520 0.915 ;
        RECT  0.310 0.305 0.410 1.310 ;
        RECT  0.065 0.305 0.310 0.495 ;
        RECT  0.185 1.210 0.310 1.310 ;
        RECT  0.065 1.210 0.185 1.460 ;
    END
END LNQD4

MACRO LNSND1
    CLASS CORE ;
    FOREIGN LNSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0464 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.680 1.770 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.310 2.575 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 0.275 3.150 1.490 ;
        RECT  2.960 0.275 3.040 0.645 ;
        RECT  2.960 1.050 3.040 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.425 0.890 1.545 ;
        RECT  0.355 1.425 0.680 1.525 ;
        RECT  0.265 0.710 0.355 1.525 ;
        RECT  0.240 0.710 0.265 1.090 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.910 0.755 1.090 ;
        RECT  0.450 0.780 0.640 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.025 1.635 3.200 1.965 ;
        RECT  1.855 1.380 2.025 1.965 ;
        RECT  0.000 1.635 1.855 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.805 0.750 2.930 0.920 ;
        RECT  2.695 0.750 2.805 1.500 ;
        RECT  2.295 1.400 2.695 1.500 ;
        RECT  2.295 0.305 2.360 0.415 ;
        RECT  2.190 0.305 2.295 1.500 ;
        RECT  1.960 0.400 2.070 1.290 ;
        RECT  1.690 0.400 1.960 0.510 ;
        RECT  1.695 1.180 1.960 1.290 ;
        RECT  1.585 1.180 1.695 1.525 ;
        RECT  1.340 1.425 1.585 1.525 ;
        RECT  1.375 0.850 1.530 1.020 ;
        RECT  1.260 0.315 1.375 1.335 ;
        RECT  1.130 1.425 1.340 1.545 ;
        RECT  0.775 0.315 1.260 0.405 ;
        RECT  0.785 1.245 1.260 1.335 ;
        RECT  1.000 1.025 1.140 1.135 ;
        RECT  0.910 0.495 1.000 1.135 ;
        RECT  0.610 0.495 0.910 0.660 ;
        RECT  0.185 0.495 0.610 0.600 ;
        RECT  0.140 0.410 0.185 0.600 ;
        RECT  0.140 1.345 0.175 1.525 ;
        RECT  0.050 0.410 0.140 1.525 ;
    END
END LNSND1

MACRO LNSND2
    CLASS CORE ;
    FOREIGN LNSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0465 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.680 1.770 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.285 2.785 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.275 3.350 1.490 ;
        RECT  3.165 0.275 3.240 0.645 ;
        RECT  3.165 1.050 3.240 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.425 0.890 1.545 ;
        RECT  0.355 1.425 0.680 1.525 ;
        RECT  0.265 0.710 0.355 1.525 ;
        RECT  0.240 0.710 0.265 1.110 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.910 0.755 1.090 ;
        RECT  0.450 0.780 0.640 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.045 1.635 3.600 1.965 ;
        RECT  1.850 1.380 2.045 1.965 ;
        RECT  0.000 1.635 1.850 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 0.750 3.130 0.920 ;
        RECT  2.910 0.750 3.020 1.500 ;
        RECT  2.310 1.400 2.910 1.500 ;
        RECT  2.185 0.255 2.310 1.500 ;
        RECT  1.940 0.400 2.030 1.290 ;
        RECT  1.660 0.400 1.940 0.510 ;
        RECT  1.695 1.180 1.940 1.290 ;
        RECT  1.585 1.180 1.695 1.525 ;
        RECT  1.340 1.425 1.585 1.525 ;
        RECT  1.375 0.850 1.530 1.020 ;
        RECT  1.260 0.315 1.375 1.335 ;
        RECT  1.130 1.425 1.340 1.545 ;
        RECT  0.770 0.315 1.260 0.405 ;
        RECT  0.775 1.245 1.260 1.335 ;
        RECT  1.000 1.025 1.140 1.135 ;
        RECT  0.910 0.495 1.000 1.135 ;
        RECT  0.610 0.495 0.910 0.660 ;
        RECT  0.185 0.495 0.610 0.600 ;
        RECT  0.140 0.410 0.185 0.600 ;
        RECT  0.140 1.345 0.175 1.525 ;
        RECT  0.050 0.410 0.140 1.525 ;
    END
END LNSND2

MACRO LNSND4
    CLASS CORE ;
    FOREIGN LNSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.700 1.950 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.310 3.715 0.695 ;
        RECT  3.450 1.110 3.715 1.290 ;
        RECT  3.150 0.310 3.450 1.290 ;
        RECT  3.025 0.310 3.150 0.695 ;
        RECT  3.025 1.110 3.150 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.310 4.750 0.690 ;
        RECT  4.650 1.110 4.750 1.490 ;
        RECT  4.350 0.310 4.650 1.490 ;
        RECT  4.025 0.310 4.350 0.690 ;
        RECT  4.025 1.110 4.350 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0781 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.425 0.880 1.545 ;
        RECT  0.355 1.425 0.670 1.525 ;
        RECT  0.265 0.710 0.355 1.525 ;
        RECT  0.230 0.710 0.265 1.110 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.910 0.755 1.090 ;
        RECT  0.450 0.780 0.640 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 5.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.025 0.310 4.250 0.690 ;
        RECT  4.025 1.110 4.250 1.490 ;
        RECT  3.550 0.310 3.715 0.695 ;
        RECT  3.550 1.110 3.715 1.290 ;
        RECT  3.025 0.310 3.050 0.695 ;
        RECT  3.025 1.110 3.050 1.290 ;
        RECT  3.915 0.800 4.160 0.910 ;
        RECT  3.825 0.800 3.915 1.505 ;
        RECT  2.675 1.400 3.825 1.505 ;
        RECT  2.780 0.600 2.890 1.200 ;
        RECT  2.675 0.600 2.780 0.690 ;
        RECT  2.675 1.110 2.780 1.200 ;
        RECT  2.565 0.310 2.675 0.690 ;
        RECT  2.565 1.110 2.675 1.505 ;
        RECT  2.475 0.800 2.670 0.910 ;
        RECT  2.365 0.345 2.475 1.505 ;
        RECT  1.765 0.345 2.365 0.455 ;
        RECT  1.715 1.395 2.365 1.505 ;
        RECT  2.145 0.700 2.255 1.285 ;
        RECT  1.520 1.180 2.145 1.285 ;
        RECT  1.525 1.395 1.715 1.525 ;
        RECT  1.320 1.425 1.525 1.525 ;
        RECT  1.410 0.315 1.520 1.285 ;
        RECT  0.770 0.315 1.410 0.405 ;
        RECT  1.375 1.180 1.410 1.285 ;
        RECT  1.260 1.180 1.375 1.335 ;
        RECT  1.110 1.425 1.320 1.545 ;
        RECT  0.775 1.245 1.260 1.335 ;
        RECT  1.000 1.025 1.120 1.135 ;
        RECT  0.910 0.495 1.000 1.135 ;
        RECT  0.610 0.495 0.910 0.660 ;
        RECT  0.185 0.495 0.610 0.600 ;
        RECT  0.140 0.395 0.185 0.600 ;
        RECT  0.140 1.345 0.175 1.525 ;
        RECT  0.050 0.395 0.140 1.525 ;
    END
END LNSND4

MACRO LNSNDD1
    CLASS CORE ;
    FOREIGN LNSNDD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.170 0.710 2.250 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.305 3.150 1.175 ;
        RECT  2.865 0.305 3.050 0.415 ;
        RECT  2.915 0.965 3.050 1.175 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.275 3.550 1.490 ;
        RECT  3.415 0.275 3.450 0.675 ;
        RECT  3.420 1.080 3.450 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.600 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.635 3.600 1.965 ;
        RECT  2.350 1.495 2.520 1.965 ;
        RECT  0.000 1.635 2.350 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.330 0.750 3.360 0.920 ;
        RECT  3.240 0.750 3.330 1.375 ;
        RECT  2.810 1.285 3.240 1.375 ;
        RECT  2.700 0.495 2.810 1.460 ;
        RECT  2.480 0.500 2.590 1.300 ;
        RECT  2.205 0.500 2.480 0.610 ;
        RECT  2.185 1.200 2.480 1.300 ;
        RECT  2.075 1.200 2.185 1.525 ;
        RECT  1.620 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.020 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.265 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.625 1.115 ;
        RECT  1.155 1.435 1.365 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.685 1.025 1.190 1.115 ;
        RECT  0.180 1.435 1.155 1.525 ;
        RECT  0.360 0.490 0.735 0.600 ;
        RECT  0.575 1.025 0.685 1.340 ;
        RECT  0.360 1.025 0.575 1.115 ;
        RECT  0.270 0.490 0.360 1.115 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNSNDD1

MACRO LNSNDD2
    CLASS CORE ;
    FOREIGN LNSNDD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.710 2.350 1.090 ;
        RECT  2.170 0.710 2.240 0.920 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.175 1.250 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.275 3.750 1.490 ;
        RECT  3.565 0.275 3.650 0.675 ;
        RECT  3.565 1.080 3.650 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 4.000 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.420 0.780 3.560 0.890 ;
        RECT  3.330 0.780 3.420 1.480 ;
        RECT  2.940 1.370 3.330 1.480 ;
        RECT  2.840 0.305 2.940 1.480 ;
        RECT  2.515 0.305 2.840 0.415 ;
        RECT  2.515 1.370 2.840 1.480 ;
        RECT  2.620 0.510 2.730 1.280 ;
        RECT  2.265 0.510 2.620 0.620 ;
        RECT  2.185 1.180 2.620 1.280 ;
        RECT  2.075 1.180 2.185 1.525 ;
        RECT  1.620 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.030 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.265 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.625 1.115 ;
        RECT  1.155 1.435 1.365 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.685 1.025 1.190 1.115 ;
        RECT  0.180 1.435 1.155 1.525 ;
        RECT  0.360 0.490 0.735 0.600 ;
        RECT  0.575 1.025 0.685 1.340 ;
        RECT  0.360 1.025 0.575 1.115 ;
        RECT  0.270 0.490 0.360 1.115 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNSNDD2

MACRO LNSNDD4
    CLASS CORE ;
    FOREIGN LNSNDD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.700 2.360 1.090 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.325 4.265 0.635 ;
        RECT  4.050 1.110 4.255 1.290 ;
        RECT  3.750 0.325 4.050 1.290 ;
        RECT  3.545 0.325 3.750 0.635 ;
        RECT  3.555 1.110 3.750 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.230 0.325 5.285 0.635 ;
        RECT  5.230 1.100 5.285 1.410 ;
        RECT  4.930 0.325 5.230 1.410 ;
        RECT  4.565 0.325 4.930 0.635 ;
        RECT  4.565 1.100 4.930 1.410 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.495 -0.165 5.600 0.165 ;
        RECT  5.385 -0.165 5.495 0.685 ;
        RECT  0.000 -0.165 5.385 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.495 1.635 5.600 1.965 ;
        RECT  5.385 1.050 5.495 1.965 ;
        RECT  0.000 1.635 5.385 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.565 0.325 4.850 0.635 ;
        RECT  4.565 1.100 4.850 1.410 ;
        RECT  4.150 0.325 4.265 0.635 ;
        RECT  4.150 1.110 4.255 1.290 ;
        RECT  3.545 0.325 3.650 0.635 ;
        RECT  3.555 1.110 3.650 1.290 ;
        RECT  4.465 0.780 4.710 0.890 ;
        RECT  4.375 0.780 4.465 1.505 ;
        RECT  3.195 1.400 4.375 1.505 ;
        RECT  3.310 0.595 3.410 1.150 ;
        RECT  3.195 0.595 3.310 0.685 ;
        RECT  3.195 1.050 3.310 1.150 ;
        RECT  3.085 0.275 3.195 0.685 ;
        RECT  3.085 1.050 3.195 1.505 ;
        RECT  2.995 0.780 3.190 0.890 ;
        RECT  2.885 0.490 2.995 1.495 ;
        RECT  2.275 0.490 2.885 0.600 ;
        RECT  1.830 1.385 2.885 1.495 ;
        RECT  2.660 0.750 2.770 1.295 ;
        RECT  2.030 1.205 2.660 1.295 ;
        RECT  1.920 0.295 2.030 1.295 ;
        RECT  1.235 0.295 1.920 0.405 ;
        RECT  1.475 1.205 1.920 1.295 ;
        RECT  1.620 1.385 1.830 1.525 ;
        RECT  1.300 1.005 1.625 1.115 ;
        RECT  1.265 1.205 1.475 1.315 ;
        RECT  1.155 1.435 1.365 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.685 1.025 1.190 1.115 ;
        RECT  0.180 1.435 1.155 1.525 ;
        RECT  0.360 0.490 0.735 0.600 ;
        RECT  0.575 1.025 0.685 1.340 ;
        RECT  0.360 1.025 0.575 1.115 ;
        RECT  0.270 0.490 0.360 1.115 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.275 0.180 0.675 ;
        RECT  0.150 1.050 0.180 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LNSNDD4

MACRO LNSNDQD1
    CLASS CORE ;
    FOREIGN LNSNDQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.170 0.710 2.250 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.150 1.490 ;
        RECT  3.015 0.275 3.050 0.675 ;
        RECT  3.015 1.080 3.050 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.165 3.200 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.200 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.920 0.750 2.960 0.920 ;
        RECT  2.820 0.305 2.920 1.495 ;
        RECT  2.465 0.305 2.820 0.415 ;
        RECT  2.485 1.385 2.820 1.495 ;
        RECT  2.600 0.510 2.710 1.290 ;
        RECT  2.215 0.510 2.600 0.620 ;
        RECT  2.165 1.190 2.600 1.290 ;
        RECT  2.055 1.190 2.165 1.525 ;
        RECT  1.600 1.415 2.055 1.525 ;
        RECT  1.920 0.750 2.010 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.245 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.605 1.115 ;
        RECT  1.135 1.435 1.345 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.685 1.025 1.190 1.115 ;
        RECT  0.180 1.435 1.135 1.525 ;
        RECT  0.360 0.490 0.735 0.600 ;
        RECT  0.575 1.025 0.685 1.340 ;
        RECT  0.360 1.025 0.575 1.115 ;
        RECT  0.270 0.490 0.360 1.115 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNSNDQD1

MACRO LNSNDQD2
    CLASS CORE ;
    FOREIGN LNSNDQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.220 0.710 2.250 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.575 3.350 1.180 ;
        RECT  3.205 0.575 3.250 0.675 ;
        RECT  3.205 1.080 3.250 1.180 ;
        RECT  3.095 0.275 3.205 0.675 ;
        RECT  3.095 1.080 3.205 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 -0.165 3.600 0.165 ;
        RECT  3.355 -0.165 3.465 0.485 ;
        RECT  0.880 -0.165 3.355 0.165 ;
        RECT  0.770 -0.165 0.880 0.355 ;
        RECT  0.000 -0.165 0.770 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 1.635 3.600 1.965 ;
        RECT  3.355 1.280 3.465 1.965 ;
        RECT  0.000 1.635 3.355 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.000 0.780 3.160 0.890 ;
        RECT  2.900 0.305 3.000 1.495 ;
        RECT  2.525 0.305 2.900 0.415 ;
        RECT  2.545 1.385 2.900 1.495 ;
        RECT  2.660 0.510 2.770 1.290 ;
        RECT  2.275 0.510 2.660 0.620 ;
        RECT  2.185 1.190 2.660 1.290 ;
        RECT  2.075 1.190 2.185 1.525 ;
        RECT  1.600 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.020 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.245 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.605 1.115 ;
        RECT  1.135 1.435 1.345 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.685 1.025 1.190 1.115 ;
        RECT  0.180 1.435 1.135 1.525 ;
        RECT  0.360 0.490 0.735 0.600 ;
        RECT  0.575 1.025 0.685 1.340 ;
        RECT  0.360 1.025 0.575 1.115 ;
        RECT  0.270 0.490 0.360 1.115 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.440 0.180 0.650 ;
        RECT  0.150 1.130 0.180 1.525 ;
        RECT  0.090 0.440 0.150 1.525 ;
        RECT  0.060 0.440 0.090 1.340 ;
    END
END LNSNDQD2

MACRO LNSNDQD4
    CLASS CORE ;
    FOREIGN LNSNDQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.350 1.090 ;
        RECT  2.220 0.710 2.250 0.920 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.325 3.750 0.635 ;
        RECT  3.650 1.100 3.750 1.410 ;
        RECT  3.350 0.325 3.650 1.410 ;
        RECT  3.015 0.325 3.350 0.635 ;
        RECT  3.015 1.100 3.350 1.410 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.920 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.050 0.890 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 4.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.015 0.325 3.250 0.635 ;
        RECT  3.015 1.100 3.250 1.410 ;
        RECT  2.905 0.780 3.160 0.890 ;
        RECT  2.805 0.305 2.905 1.495 ;
        RECT  2.515 0.305 2.805 0.415 ;
        RECT  2.535 1.385 2.805 1.495 ;
        RECT  2.585 0.510 2.695 1.290 ;
        RECT  2.265 0.510 2.585 0.620 ;
        RECT  2.185 1.190 2.585 1.290 ;
        RECT  2.075 1.190 2.185 1.525 ;
        RECT  1.600 1.415 2.075 1.525 ;
        RECT  1.920 0.750 2.020 0.920 ;
        RECT  1.820 0.295 1.920 1.315 ;
        RECT  1.235 0.295 1.820 0.405 ;
        RECT  1.245 1.205 1.820 1.315 ;
        RECT  1.300 1.005 1.605 1.115 ;
        RECT  1.135 1.435 1.345 1.545 ;
        RECT  1.190 0.505 1.300 1.115 ;
        RECT  0.685 1.025 1.190 1.115 ;
        RECT  0.180 1.435 1.135 1.525 ;
        RECT  0.360 0.490 0.735 0.600 ;
        RECT  0.575 1.025 0.685 1.340 ;
        RECT  0.360 1.025 0.575 1.115 ;
        RECT  0.270 0.490 0.360 1.115 ;
        RECT  0.240 0.750 0.270 0.920 ;
        RECT  0.150 0.275 0.180 0.675 ;
        RECT  0.150 1.050 0.180 1.525 ;
        RECT  0.060 0.275 0.150 1.525 ;
    END
END LNSNDQD4

MACRO LNSNQD1
    CLASS CORE ;
    FOREIGN LNSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0464 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.680 1.770 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.275 2.950 1.490 ;
        RECT  2.765 0.275 2.850 0.645 ;
        RECT  2.765 1.050 2.850 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.425 0.890 1.545 ;
        RECT  0.355 1.425 0.680 1.525 ;
        RECT  0.265 0.710 0.355 1.525 ;
        RECT  0.240 0.710 0.265 1.110 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.910 0.755 1.090 ;
        RECT  0.450 0.780 0.640 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.615 -0.165 3.000 0.165 ;
        RECT  2.485 -0.165 2.615 0.645 ;
        RECT  0.000 -0.165 2.485 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.615 1.635 3.000 1.965 ;
        RECT  2.485 1.050 2.615 1.965 ;
        RECT  2.025 1.635 2.485 1.965 ;
        RECT  1.855 1.380 2.025 1.965 ;
        RECT  0.000 1.635 1.855 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.335 0.760 2.740 0.910 ;
        RECT  2.190 0.270 2.335 1.500 ;
        RECT  1.960 0.400 2.070 1.290 ;
        RECT  1.690 0.400 1.960 0.510 ;
        RECT  1.695 1.180 1.960 1.290 ;
        RECT  1.585 1.180 1.695 1.525 ;
        RECT  1.340 1.425 1.585 1.525 ;
        RECT  1.375 0.850 1.530 1.020 ;
        RECT  1.260 0.315 1.375 1.335 ;
        RECT  1.130 1.425 1.340 1.545 ;
        RECT  0.775 0.315 1.260 0.405 ;
        RECT  0.785 1.245 1.260 1.335 ;
        RECT  1.000 1.025 1.140 1.135 ;
        RECT  0.910 0.495 1.000 1.135 ;
        RECT  0.610 0.495 0.910 0.660 ;
        RECT  0.185 0.495 0.610 0.600 ;
        RECT  0.140 0.410 0.185 0.600 ;
        RECT  0.140 1.345 0.175 1.525 ;
        RECT  0.050 0.410 0.140 1.525 ;
    END
END LNSNQD1

MACRO LNSNQD2
    CLASS CORE ;
    FOREIGN LNSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0465 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.680 1.770 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.540 2.950 1.185 ;
        RECT  2.830 0.540 2.840 0.645 ;
        RECT  2.830 1.050 2.840 1.185 ;
        RECT  2.710 0.275 2.830 0.645 ;
        RECT  2.710 1.050 2.830 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.425 0.890 1.545 ;
        RECT  0.355 1.425 0.680 1.525 ;
        RECT  0.265 0.710 0.355 1.525 ;
        RECT  0.240 0.710 0.265 1.110 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.910 0.755 1.090 ;
        RECT  0.450 0.780 0.640 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.090 -0.165 3.200 0.165 ;
        RECT  2.970 -0.165 3.090 0.445 ;
        RECT  2.570 -0.165 2.970 0.165 ;
        RECT  2.450 -0.165 2.570 0.645 ;
        RECT  0.000 -0.165 2.450 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.090 1.635 3.200 1.965 ;
        RECT  2.970 1.295 3.090 1.965 ;
        RECT  2.570 1.635 2.970 1.965 ;
        RECT  2.450 1.050 2.570 1.965 ;
        RECT  2.045 1.635 2.450 1.965 ;
        RECT  1.850 1.380 2.045 1.965 ;
        RECT  0.000 1.635 1.850 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.310 0.775 2.735 0.900 ;
        RECT  2.185 0.255 2.310 1.500 ;
        RECT  1.940 0.400 2.030 1.290 ;
        RECT  1.660 0.400 1.940 0.510 ;
        RECT  1.695 1.180 1.940 1.290 ;
        RECT  1.585 1.180 1.695 1.525 ;
        RECT  1.340 1.425 1.585 1.525 ;
        RECT  1.375 0.850 1.530 1.020 ;
        RECT  1.260 0.315 1.375 1.335 ;
        RECT  1.130 1.425 1.340 1.545 ;
        RECT  0.770 0.315 1.260 0.405 ;
        RECT  0.785 1.245 1.260 1.335 ;
        RECT  1.000 1.025 1.140 1.135 ;
        RECT  0.910 0.495 1.000 1.135 ;
        RECT  0.610 0.495 0.910 0.660 ;
        RECT  0.185 0.495 0.610 0.600 ;
        RECT  0.140 0.410 0.185 0.600 ;
        RECT  0.140 1.345 0.175 1.525 ;
        RECT  0.050 0.410 0.140 1.525 ;
    END
END LNSNQD2

MACRO LNSNQD4
    CLASS CORE ;
    FOREIGN LNSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0465 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.680 1.770 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.315 0.690 ;
        RECT  3.050 1.110 3.315 1.490 ;
        RECT  2.750 0.310 3.050 1.490 ;
        RECT  2.650 0.310 2.750 0.690 ;
        RECT  2.650 1.110 2.750 1.490 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0778 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.425 0.890 1.545 ;
        RECT  0.355 1.425 0.680 1.525 ;
        RECT  0.265 0.700 0.355 1.525 ;
        RECT  0.240 0.700 0.265 1.110 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.910 0.755 1.090 ;
        RECT  0.450 0.780 0.640 1.090 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.045 1.635 3.600 1.965 ;
        RECT  1.850 1.380 2.045 1.965 ;
        RECT  0.000 1.635 1.850 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 0.310 3.315 0.690 ;
        RECT  3.150 1.110 3.315 1.490 ;
        RECT  2.310 0.800 2.640 0.900 ;
        RECT  2.185 0.255 2.310 1.525 ;
        RECT  1.920 0.400 2.050 1.290 ;
        RECT  1.660 0.400 1.920 0.510 ;
        RECT  1.695 1.180 1.920 1.290 ;
        RECT  1.585 1.180 1.695 1.525 ;
        RECT  1.340 1.425 1.585 1.525 ;
        RECT  1.375 0.850 1.530 1.020 ;
        RECT  1.260 0.315 1.375 1.335 ;
        RECT  1.130 1.425 1.340 1.545 ;
        RECT  0.770 0.315 1.260 0.405 ;
        RECT  0.785 1.245 1.260 1.335 ;
        RECT  1.000 1.025 1.140 1.135 ;
        RECT  0.910 0.495 1.000 1.135 ;
        RECT  0.610 0.495 0.910 0.660 ;
        RECT  0.185 0.495 0.610 0.590 ;
        RECT  0.140 0.395 0.185 0.590 ;
        RECT  0.140 1.345 0.175 1.525 ;
        RECT  0.050 0.395 0.140 1.525 ;
    END
END LNSNQD4

MACRO LVLHLD1
    CLASS CORE ;
    FOREIGN LVLHLD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.310 0.750 1.490 ;
        RECT  0.610 0.310 0.650 0.520 ;
        RECT  0.610 1.060 0.650 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.180 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 -0.165 0.800 0.165 ;
        RECT  0.315 -0.165 0.500 0.420 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.635 0.800 1.965 ;
        RECT  0.315 1.380 0.495 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.475 0.730 0.555 0.940 ;
        RECT  0.375 0.510 0.475 1.290 ;
        RECT  0.200 0.510 0.375 0.600 ;
        RECT  0.200 1.200 0.375 1.290 ;
        RECT  0.090 0.280 0.200 0.600 ;
        RECT  0.090 1.200 0.200 1.490 ;
    END
END LVLHLD1

MACRO LVLHLD2
    CLASS CORE ;
    FOREIGN LVLHLD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.275 0.760 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.195 0.940 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.165 1.200 0.165 ;
        RECT  0.905 -0.165 1.015 0.695 ;
        RECT  0.500 -0.165 0.905 0.165 ;
        RECT  0.330 -0.165 0.500 0.390 ;
        RECT  0.000 -0.165 0.330 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 1.635 1.200 1.965 ;
        RECT  0.905 1.040 1.015 1.965 ;
        RECT  0.500 1.635 0.905 1.965 ;
        RECT  0.330 1.410 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.420 0.500 0.530 1.300 ;
        RECT  0.185 0.500 0.420 0.600 ;
        RECT  0.185 1.200 0.420 1.300 ;
        RECT  0.075 0.390 0.185 0.600 ;
        RECT  0.075 1.200 0.185 1.425 ;
    END
END LVLHLD2

MACRO LVLHLD4
    CLASS CORE ;
    FOREIGN LVLHLD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.310 1.450 1.490 ;
        RECT  0.845 0.310 1.150 0.690 ;
        RECT  0.845 1.110 1.150 1.490 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.785 0.505 0.890 ;
        RECT  0.050 0.700 0.155 1.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 -0.165 1.800 0.165 ;
        RECT  1.605 -0.165 1.715 0.690 ;
        RECT  0.195 -0.165 1.605 0.165 ;
        RECT  0.085 -0.165 0.195 0.525 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.635 1.800 1.965 ;
        RECT  1.605 1.110 1.715 1.965 ;
        RECT  0.195 1.635 1.605 1.965 ;
        RECT  0.085 1.260 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.845 0.310 1.050 0.690 ;
        RECT  0.845 1.110 1.050 1.490 ;
        RECT  0.730 0.780 0.925 0.890 ;
        RECT  0.630 0.585 0.730 1.150 ;
        RECT  0.455 0.585 0.630 0.695 ;
        RECT  0.455 1.040 0.630 1.150 ;
        RECT  0.345 0.275 0.455 0.695 ;
        RECT  0.345 1.040 0.455 1.470 ;
    END
END LVLHLD4

MACRO LVLHLD8
    CLASS CORE ;
    FOREIGN LVLHLD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.325 2.850 0.690 ;
        RECT  2.250 1.110 2.845 1.475 ;
        RECT  1.750 0.325 2.250 1.475 ;
        RECT  1.100 0.325 1.750 0.690 ;
        RECT  1.100 1.110 1.750 1.475 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.780 0.760 0.890 ;
        RECT  0.250 0.700 0.350 1.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.165 3.200 0.165 ;
        RECT  2.960 -0.165 3.070 0.695 ;
        RECT  0.000 -0.165 2.960 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 1.635 3.200 1.965 ;
        RECT  2.960 1.040 3.070 1.965 ;
        RECT  0.990 1.635 2.960 1.965 ;
        RECT  0.880 1.260 0.990 1.965 ;
        RECT  0.000 1.635 0.880 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.325 2.850 0.690 ;
        RECT  2.350 1.110 2.845 1.475 ;
        RECT  1.100 0.325 1.650 0.690 ;
        RECT  1.100 1.110 1.650 1.475 ;
        RECT  2.495 0.800 2.925 0.910 ;
        RECT  0.990 0.800 1.460 0.910 ;
        RECT  0.890 0.580 0.990 1.150 ;
        RECT  0.730 0.580 0.890 0.690 ;
        RECT  0.730 1.040 0.890 1.150 ;
        RECT  0.620 0.295 0.730 0.690 ;
        RECT  0.620 1.040 0.730 1.470 ;
        RECT  0.050 0.385 0.620 0.495 ;
        RECT  0.050 1.360 0.620 1.470 ;
    END
END LVLHLD8

MACRO LVLLHCD1
    CLASS CORE ;
    FOREIGN LVLLHCD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.1710 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 2.900 2.550 3.000 ;
        RECT  2.050 2.310 2.190 3.290 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 2.600 3.150 3.090 ;
        RECT  2.700 2.600 3.050 2.710 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.1248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.265 1.635 3.600 1.965 ;
        RECT  3.155 1.635 3.265 2.275 ;
        RECT  2.745 1.635 3.155 1.965 ;
        RECT  2.635 1.635 2.745 2.275 ;
        RECT  0.000 1.635 2.635 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 3.600 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.600 0.165 ;
        RECT  2.740 3.435 3.600 3.765 ;
        RECT  2.640 2.845 2.740 3.765 ;
        RECT  1.935 3.435 2.640 3.765 ;
        RECT  1.825 2.910 1.935 3.765 ;
        RECT  0.000 3.435 1.825 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.415 2.110 3.525 2.490 ;
        RECT  3.005 2.400 3.415 2.490 ;
        RECT  2.895 2.110 3.005 2.490 ;
        RECT  2.485 2.400 2.895 2.490 ;
        RECT  2.410 1.415 2.545 1.525 ;
        RECT  2.375 2.110 2.485 2.490 ;
        RECT  2.300 1.000 2.410 1.525 ;
        RECT  0.295 2.110 2.375 2.220 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.850 2.530 1.960 2.790 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.715 2.680 1.850 2.790 ;
        RECT  0.940 2.345 1.785 2.455 ;
        RECT  1.605 2.680 1.715 3.290 ;
        RECT  1.060 2.770 1.605 2.870 ;
        RECT  0.185 3.200 1.605 3.290 ;
        RECT  0.940 2.995 1.265 3.105 ;
        RECT  0.850 2.345 0.940 3.105 ;
        RECT  0.755 2.725 0.850 2.915 ;
        RECT  0.185 2.345 0.740 2.455 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.075 2.110 0.185 3.290 ;
    END
END LVLLHCD1

MACRO LVLLHCD2
    CLASS CORE ;
    FOREIGN LVLLHCD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.2360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 2.820 3.185 2.920 ;
        RECT  2.420 2.310 2.550 3.290 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.1400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 2.600 3.550 3.090 ;
        RECT  3.110 2.600 3.450 2.710 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.1248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.655 1.635 4.000 1.965 ;
        RECT  3.545 1.635 3.655 2.275 ;
        RECT  3.135 1.635 3.545 1.965 ;
        RECT  3.025 1.635 3.135 2.275 ;
        RECT  0.000 1.635 3.025 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 4.000 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.000 0.165 ;
        RECT  2.785 3.435 4.000 3.765 ;
        RECT  2.675 3.095 2.785 3.765 ;
        RECT  2.265 3.435 2.675 3.765 ;
        RECT  2.155 2.910 2.265 3.765 ;
        RECT  0.000 3.435 2.155 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.805 2.110 3.915 2.490 ;
        RECT  3.395 2.400 3.805 2.490 ;
        RECT  3.285 2.110 3.395 2.490 ;
        RECT  2.830 2.400 3.285 2.490 ;
        RECT  2.720 2.110 2.830 2.490 ;
        RECT  2.265 2.110 2.720 2.220 ;
        RECT  2.410 1.415 2.565 1.525 ;
        RECT  2.300 1.000 2.410 1.525 ;
        RECT  2.060 2.600 2.310 2.700 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  2.155 2.110 2.265 2.490 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  1.225 2.110 2.155 2.220 ;
        RECT  1.960 2.600 2.060 3.290 ;
        RECT  1.440 2.345 2.045 2.455 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.595 2.770 1.960 2.870 ;
        RECT  0.405 3.200 1.960 3.290 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.440 2.995 1.850 3.105 ;
        RECT  1.335 2.345 1.440 3.105 ;
        RECT  1.115 2.110 1.225 2.455 ;
        RECT  0.185 2.110 1.115 2.220 ;
        RECT  0.405 2.345 1.005 2.455 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.295 2.345 0.405 3.290 ;
        RECT  0.075 2.110 0.185 2.490 ;
    END
END LVLLHCD2

MACRO LVLLHCD4
    CLASS CORE ;
    FOREIGN LVLLHCD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.4470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 2.910 2.810 3.290 ;
        RECT  2.050 2.310 2.305 2.490 ;
        RECT  1.750 2.310 2.050 3.290 ;
        RECT  1.595 2.310 1.750 2.490 ;
        RECT  1.595 2.910 1.750 3.290 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.2206 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 2.910 3.970 3.290 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.1248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.045 1.635 4.200 1.965 ;
        RECT  3.935 1.635 4.045 2.490 ;
        RECT  0.000 1.635 3.935 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 4.200 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.200 0.165 ;
        RECT  0.000 3.435 4.200 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.150 2.910 2.810 3.290 ;
        RECT  2.150 2.310 2.305 2.490 ;
        RECT  1.595 2.310 1.650 2.490 ;
        RECT  1.595 2.910 1.650 3.290 ;
        RECT  3.675 2.110 3.785 2.735 ;
        RECT  3.285 2.645 3.675 2.735 ;
        RECT  3.175 2.110 3.285 2.735 ;
        RECT  2.785 2.645 3.175 2.735 ;
        RECT  2.675 2.110 2.785 2.735 ;
        RECT  2.525 2.110 2.675 2.220 ;
        RECT  2.410 1.415 2.565 1.525 ;
        RECT  2.415 2.110 2.525 2.490 ;
        RECT  1.485 2.110 2.415 2.220 ;
        RECT  2.300 1.000 2.410 1.525 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.485 2.600 1.640 2.700 ;
        RECT  1.375 2.110 1.485 2.490 ;
        RECT  1.375 2.600 1.485 3.290 ;
        RECT  0.295 2.110 1.375 2.220 ;
        RECT  1.060 2.770 1.375 2.870 ;
        RECT  0.185 3.200 1.375 3.290 ;
        RECT  0.940 2.345 1.265 2.455 ;
        RECT  0.940 2.995 1.265 3.105 ;
        RECT  0.850 2.345 0.940 3.105 ;
        RECT  0.755 2.725 0.850 2.915 ;
        RECT  0.185 2.345 0.740 2.455 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.075 2.110 0.185 3.290 ;
    END
END LVLLHCD4

MACRO LVLLHCD8
    CLASS CORE ;
    FOREIGN LVLLHCD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.8320 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 2.910 4.565 3.275 ;
        RECT  3.450 2.350 4.125 2.490 ;
        RECT  2.950 2.350 3.450 3.275 ;
        RECT  2.375 2.350 2.950 2.490 ;
        RECT  2.375 2.910 2.950 3.275 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.4391 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 2.845 6.760 3.290 ;
        RECT  5.150 3.200 6.650 3.290 ;
        RECT  5.020 2.845 5.150 3.290 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.1482 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.845 1.635 7.000 1.965 ;
        RECT  6.735 1.635 6.845 2.490 ;
        RECT  6.325 1.635 6.735 1.965 ;
        RECT  6.215 1.635 6.325 2.490 ;
        RECT  5.805 1.635 6.215 1.965 ;
        RECT  5.695 1.635 5.805 2.490 ;
        RECT  5.285 1.635 5.695 1.965 ;
        RECT  5.175 1.635 5.285 2.490 ;
        RECT  4.765 1.635 5.175 1.965 ;
        RECT  4.655 1.635 4.765 2.490 ;
        RECT  0.000 1.635 4.655 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 7.000 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 7.000 0.165 ;
        RECT  4.785 3.435 7.000 3.765 ;
        RECT  4.675 2.910 4.785 3.765 ;
        RECT  2.265 3.435 4.675 3.765 ;
        RECT  2.155 2.910 2.265 3.765 ;
        RECT  0.000 3.435 2.155 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.550 2.910 4.565 3.275 ;
        RECT  3.550 2.350 4.125 2.490 ;
        RECT  2.375 2.350 2.850 2.490 ;
        RECT  2.375 2.910 2.850 3.275 ;
        RECT  6.475 2.110 6.585 2.735 ;
        RECT  6.065 2.645 6.475 2.735 ;
        RECT  5.955 2.110 6.065 2.735 ;
        RECT  5.545 2.645 5.955 2.735 ;
        RECT  5.435 2.110 5.545 2.735 ;
        RECT  5.025 2.645 5.435 2.735 ;
        RECT  4.915 2.110 5.025 2.735 ;
        RECT  4.505 2.645 4.915 2.735 ;
        RECT  4.395 2.100 4.505 2.735 ;
        RECT  2.265 2.100 4.395 2.190 ;
        RECT  3.750 2.600 4.190 2.700 ;
        RECT  2.060 2.600 2.750 2.700 ;
        RECT  2.410 1.415 2.565 1.525 ;
        RECT  2.300 1.000 2.410 1.525 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  2.155 2.100 2.265 2.490 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  1.225 2.110 2.155 2.220 ;
        RECT  1.960 2.600 2.060 3.290 ;
        RECT  1.440 2.345 2.045 2.455 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.595 2.770 1.960 2.870 ;
        RECT  0.405 3.200 1.960 3.290 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.440 2.995 1.850 3.105 ;
        RECT  1.335 2.345 1.440 3.105 ;
        RECT  1.115 2.110 1.225 2.455 ;
        RECT  0.185 2.110 1.115 2.220 ;
        RECT  0.405 2.345 1.005 2.455 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.295 2.345 0.405 3.290 ;
        RECT  0.075 2.110 0.185 2.490 ;
    END
END LVLLHCD8

MACRO LVLLHD1
    CLASS CORE ;
    FOREIGN LVLLHD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.1580 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 2.110 2.350 3.290 ;
        RECT  2.150 2.110 2.240 2.490 ;
        RECT  2.150 2.910 2.240 3.290 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.635 2.600 1.965 ;
        RECT  2.300 1.000 2.410 1.965 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  1.995 1.635 2.300 1.965 ;
        RECT  1.885 1.635 1.995 2.290 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.485 1.635 1.885 1.965 ;
        RECT  1.375 1.635 1.485 2.290 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.855 1.635 0.965 2.290 ;
        RECT  0.445 1.635 0.855 1.965 ;
        RECT  0.335 1.635 0.445 2.290 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 2.600 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.600 0.165 ;
        RECT  1.995 3.435 2.600 3.765 ;
        RECT  1.885 2.910 1.995 3.765 ;
        RECT  0.000 3.435 1.885 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  1.930 2.530 2.040 2.790 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.775 2.680 1.930 2.790 ;
        RECT  1.665 2.680 1.775 3.290 ;
        RECT  1.635 2.110 1.745 2.490 ;
        RECT  1.060 2.770 1.665 2.870 ;
        RECT  0.185 3.200 1.665 3.290 ;
        RECT  1.225 2.380 1.635 2.490 ;
        RECT  0.940 2.995 1.265 3.105 ;
        RECT  1.115 2.110 1.225 2.490 ;
        RECT  0.940 2.380 1.115 2.490 ;
        RECT  0.850 2.380 0.940 3.105 ;
        RECT  0.755 2.725 0.850 2.915 ;
        RECT  0.595 2.110 0.705 2.490 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.185 2.380 0.595 2.490 ;
        RECT  0.075 2.110 0.185 3.290 ;
    END
END LVLLHD1

MACRO LVLLHD2
    CLASS CORE ;
    FOREIGN LVLLHD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 2.110 1.755 3.290 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.635 2.600 1.965 ;
        RECT  2.300 1.000 2.410 1.965 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  2.005 1.635 2.300 1.965 ;
        RECT  1.895 1.635 2.005 2.490 ;
        RECT  1.485 1.635 1.895 1.965 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.375 1.635 1.485 2.290 ;
        RECT  0.760 1.635 1.375 1.965 ;
        RECT  0.760 2.145 1.005 2.255 ;
        RECT  0.640 1.635 0.760 2.255 ;
        RECT  0.000 1.635 0.640 1.965 ;
        RECT  0.295 2.145 0.640 2.255 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 2.600 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.600 0.165 ;
        RECT  2.005 3.435 2.600 3.765 ;
        RECT  1.895 2.910 2.005 3.765 ;
        RECT  0.000 3.435 1.895 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.435 2.530 1.555 3.290 ;
        RECT  1.060 2.770 1.435 2.870 ;
        RECT  0.185 3.200 1.435 3.290 ;
        RECT  0.940 2.995 1.265 3.105 ;
        RECT  1.115 2.110 1.225 2.490 ;
        RECT  0.940 2.380 1.115 2.490 ;
        RECT  0.850 2.380 0.940 3.105 ;
        RECT  0.755 2.725 0.850 2.915 ;
        RECT  0.185 2.345 0.740 2.455 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.075 2.110 0.185 3.290 ;
    END
END LVLLHD2

MACRO LVLLHD4
    CLASS CORE ;
    FOREIGN LVLLHD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 2.110 2.305 2.490 ;
        RECT  2.050 2.910 2.305 3.290 ;
        RECT  1.750 2.110 2.050 3.290 ;
        RECT  1.595 2.110 1.750 2.490 ;
        RECT  1.595 2.910 1.750 3.290 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.525 1.635 2.600 1.965 ;
        RECT  2.415 1.635 2.525 2.490 ;
        RECT  2.410 1.635 2.415 1.965 ;
        RECT  2.300 1.000 2.410 1.965 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  1.485 1.635 2.300 1.965 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.375 1.635 1.485 2.490 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.855 1.635 0.965 2.290 ;
        RECT  0.445 1.635 0.855 1.965 ;
        RECT  0.335 1.635 0.445 2.290 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 2.600 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.600 0.165 ;
        RECT  2.525 3.435 2.600 3.765 ;
        RECT  2.415 2.910 2.525 3.765 ;
        RECT  0.000 3.435 2.415 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.150 2.110 2.305 2.490 ;
        RECT  2.150 2.910 2.305 3.290 ;
        RECT  1.595 2.110 1.650 2.490 ;
        RECT  1.595 2.910 1.650 3.290 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.485 2.600 1.640 2.700 ;
        RECT  1.375 2.600 1.485 3.290 ;
        RECT  1.060 2.770 1.375 2.870 ;
        RECT  0.185 3.200 1.375 3.290 ;
        RECT  0.950 2.995 1.265 3.105 ;
        RECT  1.115 2.110 1.225 2.490 ;
        RECT  0.950 2.380 1.115 2.490 ;
        RECT  0.850 2.380 0.950 3.105 ;
        RECT  0.755 2.725 0.850 2.915 ;
        RECT  0.595 2.110 0.705 2.490 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.185 2.380 0.595 2.490 ;
        RECT  0.075 2.110 0.185 3.290 ;
    END
END LVLLHD4

MACRO LVLLHD8
    CLASS CORE ;
    FOREIGN LVLLHD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 2.125 4.085 2.490 ;
        RECT  3.450 2.910 4.085 3.275 ;
        RECT  2.950 2.125 3.450 3.275 ;
        RECT  2.365 2.125 2.950 2.490 ;
        RECT  2.365 2.910 2.950 3.275 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1482 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 2.150 0.910 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.305 1.635 4.400 1.965 ;
        RECT  4.195 1.635 4.305 2.490 ;
        RECT  2.410 1.635 4.195 1.965 ;
        RECT  2.300 1.000 2.410 1.965 ;
        RECT  1.890 1.000 2.300 1.110 ;
        RECT  2.255 1.635 2.300 1.965 ;
        RECT  2.145 1.635 2.255 2.490 ;
        RECT  1.745 1.635 2.145 1.965 ;
        RECT  1.780 1.000 1.890 1.290 ;
        RECT  1.635 1.635 1.745 2.290 ;
        RECT  1.225 1.635 1.635 1.965 ;
        RECT  1.115 1.635 1.225 2.490 ;
        RECT  0.705 1.635 1.115 1.965 ;
        RECT  0.595 1.635 0.705 2.290 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.635 0.185 2.490 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.310 4.400 0.600 ;
        RECT  0.950 1.110 1.440 1.290 ;
        RECT  0.760 0.310 0.950 1.290 ;
        RECT  0.430 0.310 0.760 0.600 ;
        RECT  0.240 0.310 0.430 1.290 ;
        RECT  0.000 0.310 0.240 0.600 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 4.400 0.165 ;
        RECT  4.305 3.435 4.400 3.765 ;
        RECT  4.195 2.910 4.305 3.765 ;
        RECT  2.255 3.435 4.195 3.765 ;
        RECT  2.145 2.910 2.255 3.765 ;
        RECT  0.000 3.435 2.145 3.765 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.550 2.125 4.085 2.490 ;
        RECT  3.550 2.910 4.085 3.275 ;
        RECT  2.365 2.125 2.850 2.490 ;
        RECT  2.365 2.910 2.850 3.275 ;
        RECT  3.710 2.600 4.150 2.700 ;
        RECT  2.050 2.600 2.740 2.700 ;
        RECT  2.000 1.200 2.190 1.525 ;
        RECT  1.960 2.600 2.050 3.290 ;
        RECT  1.895 2.110 2.005 2.490 ;
        RECT  0.650 1.415 2.000 1.525 ;
        RECT  1.585 2.770 1.960 2.870 ;
        RECT  0.445 3.200 1.960 3.290 ;
        RECT  1.485 2.380 1.895 2.490 ;
        RECT  1.445 2.995 1.850 3.105 ;
        RECT  1.445 2.110 1.485 2.490 ;
        RECT  1.335 2.110 1.445 3.105 ;
        RECT  0.855 2.110 0.965 2.490 ;
        RECT  0.445 2.380 0.855 2.490 ;
        RECT  0.540 1.110 0.650 1.525 ;
        RECT  0.335 2.110 0.445 3.290 ;
    END
END LVLLHD8

MACRO MAOI222D0
    CLASS CORE ;
    FOREIGN MAOI222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.495 1.550 1.300 ;
        RECT  1.055 0.495 1.450 0.600 ;
        RECT  0.195 1.210 1.450 1.300 ;
        RECT  0.150 0.490 0.265 0.600 ;
        RECT  0.150 1.210 0.195 1.495 ;
        RECT  0.050 0.490 0.150 1.495 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.100 ;
        RECT  0.690 1.010 1.245 1.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.710 1.155 0.900 ;
        RECT  0.600 0.810 1.020 0.900 ;
        RECT  0.550 0.710 0.600 0.900 ;
        RECT  0.450 0.710 0.550 1.090 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.355 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.645 -0.165 1.600 0.165 ;
        RECT  0.645 0.495 0.745 0.600 ;
        RECT  0.535 -0.165 0.645 0.600 ;
        RECT  0.000 -0.165 0.535 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.635 1.600 1.965 ;
        RECT  0.595 1.405 0.705 1.965 ;
        RECT  0.515 1.405 0.595 1.515 ;
        RECT  0.000 1.635 0.595 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.275 1.540 0.385 ;
        RECT  0.795 1.410 1.540 1.520 ;
        RECT  0.845 0.275 0.955 0.645 ;
    END
END MAOI222D0

MACRO MAOI222D1
    CLASS CORE ;
    FOREIGN MAOI222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2960 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.495 1.550 1.300 ;
        RECT  1.075 0.495 1.445 0.585 ;
        RECT  0.195 1.210 1.445 1.300 ;
        RECT  0.150 0.295 0.195 0.600 ;
        RECT  0.150 1.210 0.195 1.500 ;
        RECT  0.050 0.295 0.150 1.500 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0399 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.100 ;
        RECT  0.900 1.010 1.245 1.100 ;
        RECT  0.730 0.875 0.900 1.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0809 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.695 1.155 0.900 ;
        RECT  0.620 0.695 1.010 0.785 ;
        RECT  0.570 0.695 0.620 0.920 ;
        RECT  0.445 0.695 0.570 1.090 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1016 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.355 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 -0.165 1.600 0.165 ;
        RECT  0.530 0.495 0.715 0.585 ;
        RECT  0.440 -0.165 0.530 0.585 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 1.635 1.600 1.965 ;
        RECT  0.535 1.410 0.725 1.965 ;
        RECT  0.000 1.635 0.535 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 0.295 1.525 0.385 ;
        RECT  0.815 1.410 1.525 1.500 ;
        RECT  0.895 0.295 0.985 0.585 ;
        RECT  0.815 0.480 0.895 0.585 ;
    END
END MAOI222D1

MACRO MAOI222D2
    CLASS CORE ;
    FOREIGN MAOI222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.545 2.355 1.195 ;
        RECT  2.245 0.275 2.280 1.490 ;
        RECT  2.135 0.275 2.245 0.675 ;
        RECT  2.135 1.045 2.245 1.490 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0399 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.100 ;
        RECT  0.900 1.010 1.245 1.100 ;
        RECT  0.730 0.875 0.900 1.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0809 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.695 1.155 0.900 ;
        RECT  0.620 0.695 1.010 0.785 ;
        RECT  0.570 0.695 0.620 0.920 ;
        RECT  0.445 0.695 0.570 1.090 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1016 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.355 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.535 -0.165 2.600 0.165 ;
        RECT  2.405 -0.165 2.535 0.455 ;
        RECT  2.010 -0.165 2.405 0.165 ;
        RECT  1.880 -0.165 2.010 0.455 ;
        RECT  0.530 -0.165 1.880 0.165 ;
        RECT  0.530 0.495 0.715 0.585 ;
        RECT  0.440 -0.165 0.530 0.585 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.535 1.635 2.600 1.965 ;
        RECT  2.405 1.345 2.535 1.965 ;
        RECT  2.005 1.635 2.405 1.965 ;
        RECT  1.875 1.345 2.005 1.965 ;
        RECT  0.715 1.635 1.875 1.965 ;
        RECT  0.545 1.410 0.715 1.965 ;
        RECT  0.000 1.635 0.545 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.990 0.770 2.120 0.900 ;
        RECT  1.900 0.545 1.990 1.195 ;
        RECT  1.735 0.545 1.900 0.675 ;
        RECT  1.735 1.045 1.900 1.195 ;
        RECT  1.535 0.790 1.780 0.880 ;
        RECT  1.635 0.275 1.735 0.675 ;
        RECT  1.635 1.045 1.735 1.490 ;
        RECT  1.445 0.495 1.535 1.300 ;
        RECT  0.985 0.295 1.515 0.385 ;
        RECT  1.075 0.495 1.445 0.585 ;
        RECT  0.195 1.210 1.445 1.300 ;
        RECT  0.895 0.295 0.985 0.585 ;
        RECT  0.815 0.480 0.895 0.585 ;
        RECT  0.150 0.295 0.195 0.600 ;
        RECT  0.150 1.210 0.195 1.500 ;
        RECT  0.060 0.295 0.150 1.500 ;
        RECT  0.805 1.410 1.515 1.500 ;
    END
END MAOI222D2

MACRO MAOI222D4
    CLASS CORE ;
    FOREIGN MAOI222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.310 2.895 0.690 ;
        RECT  2.650 1.110 2.895 1.490 ;
        RECT  2.350 0.310 2.650 1.490 ;
        RECT  2.115 0.310 2.350 0.690 ;
        RECT  2.115 1.110 2.350 1.490 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0399 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.350 1.100 ;
        RECT  0.900 1.010 1.245 1.100 ;
        RECT  0.730 0.875 0.900 1.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0809 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.695 1.155 0.900 ;
        RECT  0.620 0.695 1.010 0.785 ;
        RECT  0.570 0.695 0.620 0.920 ;
        RECT  0.445 0.695 0.570 1.090 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1016 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.355 1.090 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.125 -0.165 3.200 0.165 ;
        RECT  3.005 -0.165 3.125 0.690 ;
        RECT  2.005 -0.165 3.005 0.165 ;
        RECT  1.885 -0.165 2.005 0.465 ;
        RECT  0.530 -0.165 1.885 0.165 ;
        RECT  0.530 0.495 0.715 0.585 ;
        RECT  0.440 -0.165 0.530 0.585 ;
        RECT  0.000 -0.165 0.440 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.125 1.635 3.200 1.965 ;
        RECT  3.005 1.110 3.125 1.965 ;
        RECT  2.005 1.635 3.005 1.965 ;
        RECT  1.885 1.335 2.005 1.965 ;
        RECT  0.715 1.635 1.885 1.965 ;
        RECT  0.545 1.410 0.715 1.965 ;
        RECT  0.000 1.635 0.545 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 0.310 2.895 0.690 ;
        RECT  2.750 1.110 2.895 1.490 ;
        RECT  2.115 0.310 2.250 0.690 ;
        RECT  2.115 1.110 2.250 1.490 ;
        RECT  1.990 0.800 2.130 0.900 ;
        RECT  1.900 0.555 1.990 1.245 ;
        RECT  1.735 0.555 1.900 0.690 ;
        RECT  1.735 1.110 1.900 1.245 ;
        RECT  1.530 0.800 1.780 0.900 ;
        RECT  1.635 0.310 1.735 0.690 ;
        RECT  1.635 1.110 1.735 1.490 ;
        RECT  1.440 0.495 1.530 1.300 ;
        RECT  0.985 0.295 1.515 0.385 ;
        RECT  1.075 0.495 1.440 0.585 ;
        RECT  0.195 1.210 1.440 1.300 ;
        RECT  0.895 0.295 0.985 0.585 ;
        RECT  0.815 0.480 0.895 0.585 ;
        RECT  0.150 0.295 0.195 0.600 ;
        RECT  0.150 1.210 0.195 1.500 ;
        RECT  0.060 0.295 0.150 1.500 ;
        RECT  0.805 1.410 1.515 1.500 ;
    END
END MAOI222D4

MACRO MAOI22D0
    CLASS CORE ;
    FOREIGN MAOI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1040 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.290 ;
        RECT  0.965 0.510 1.450 0.600 ;
        RECT  1.040 1.200 1.450 1.290 ;
        RECT  0.850 0.285 0.965 0.600 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.880 0.565 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.980 0.880 1.050 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 -0.165 1.600 0.165 ;
        RECT  1.395 -0.165 1.505 0.400 ;
        RECT  0.705 -0.165 1.395 0.165 ;
        RECT  1.295 0.290 1.395 0.400 ;
        RECT  0.595 -0.165 0.705 0.465 ;
        RECT  0.185 -0.165 0.595 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.695 1.635 1.600 1.965 ;
        RECT  0.575 1.400 0.695 1.965 ;
        RECT  0.475 1.400 0.575 1.510 ;
        RECT  0.000 1.635 0.575 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.905 1.400 1.535 1.510 ;
        RECT  0.790 1.320 0.905 1.510 ;
        RECT  0.745 0.930 0.870 1.040 ;
        RECT  0.655 0.575 0.745 1.040 ;
        RECT  0.445 0.575 0.655 0.685 ;
        RECT  0.360 0.285 0.445 0.685 ;
        RECT  0.335 0.285 0.360 1.290 ;
        RECT  0.270 0.575 0.335 1.290 ;
        RECT  0.185 1.200 0.270 1.290 ;
        RECT  0.075 1.200 0.185 1.520 ;
    END
END MAOI22D0

MACRO MAOI22D1
    CLASS CORE ;
    FOREIGN MAOI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.505 1.550 1.295 ;
        RECT  0.960 0.505 1.450 0.595 ;
        RECT  1.035 1.205 1.450 1.295 ;
        RECT  0.850 0.290 0.960 0.595 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.565 1.120 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.090 ;
        RECT  0.970 0.710 1.045 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 1.600 0.165 ;
        RECT  0.555 -0.165 0.745 0.415 ;
        RECT  0.180 -0.165 0.555 0.165 ;
        RECT  0.065 -0.165 0.180 0.530 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.635 1.600 1.965 ;
        RECT  0.520 1.260 0.650 1.965 ;
        RECT  0.000 1.635 0.520 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.905 1.405 1.505 1.525 ;
        RECT  0.790 1.205 0.905 1.525 ;
        RECT  0.745 0.750 0.810 0.930 ;
        RECT  0.655 0.505 0.745 0.930 ;
        RECT  0.360 0.505 0.655 0.595 ;
        RECT  0.270 0.505 0.360 1.315 ;
        RECT  0.195 1.200 0.270 1.315 ;
        RECT  0.065 1.200 0.195 1.515 ;
    END
END MAOI22D1

MACRO MAOI22D2
    CLASS CORE ;
    FOREIGN MAOI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.955 0.275 2.015 0.670 ;
        RECT  1.955 1.045 2.015 1.490 ;
        RECT  1.900 0.275 1.955 1.490 ;
        RECT  1.845 0.510 1.900 1.195 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.090 ;
        RECT  0.970 0.710 1.045 0.925 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.555 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 -0.165 2.400 0.165 ;
        RECT  2.155 -0.165 2.275 0.670 ;
        RECT  1.785 -0.165 2.155 0.165 ;
        RECT  1.615 -0.165 1.785 0.400 ;
        RECT  0.680 -0.165 1.615 0.165 ;
        RECT  0.490 -0.165 0.680 0.400 ;
        RECT  0.000 -0.165 0.490 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 1.635 2.400 1.965 ;
        RECT  2.160 1.045 2.275 1.965 ;
        RECT  1.785 1.635 2.160 1.965 ;
        RECT  1.615 1.380 1.785 1.965 ;
        RECT  1.485 1.635 1.615 1.965 ;
        RECT  1.305 1.380 1.485 1.965 ;
        RECT  0.745 1.635 1.305 1.965 ;
        RECT  0.555 1.380 0.745 1.965 ;
        RECT  0.195 1.635 0.555 1.965 ;
        RECT  0.070 1.355 0.195 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.535 0.490 1.675 1.290 ;
        RECT  1.035 0.490 1.535 0.590 ;
        RECT  0.960 1.200 1.535 1.290 ;
        RECT  0.905 0.275 1.490 0.400 ;
        RECT  0.955 1.200 0.960 1.475 ;
        RECT  0.850 1.045 0.955 1.475 ;
        RECT  0.790 0.275 0.905 0.590 ;
        RECT  0.745 0.745 0.810 0.925 ;
        RECT  0.655 0.745 0.745 1.290 ;
        RECT  0.360 1.200 0.655 1.290 ;
        RECT  0.270 0.510 0.360 1.290 ;
        RECT  0.185 0.510 0.270 0.600 ;
        RECT  0.075 0.325 0.185 0.600 ;
    END
END MAOI22D2

MACRO MAOI22D4
    CLASS CORE ;
    FOREIGN MAOI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.310 2.505 0.690 ;
        RECT  2.250 1.110 2.505 1.490 ;
        RECT  1.950 0.310 2.250 1.490 ;
        RECT  1.795 0.310 1.950 0.690 ;
        RECT  1.795 1.110 1.950 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.370 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.150 1.090 ;
        RECT  0.970 0.710 1.045 0.925 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.565 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.735 -0.165 2.800 0.165 ;
        RECT  2.615 -0.165 2.735 0.700 ;
        RECT  0.655 -0.165 2.615 0.165 ;
        RECT  0.515 -0.165 0.655 0.565 ;
        RECT  0.000 -0.165 0.515 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.735 1.635 2.800 1.965 ;
        RECT  2.615 1.090 2.735 1.965 ;
        RECT  1.630 1.635 2.615 1.965 ;
        RECT  1.420 1.380 1.630 1.965 ;
        RECT  0.740 1.635 1.420 1.965 ;
        RECT  0.555 1.380 0.740 1.965 ;
        RECT  0.195 1.635 0.555 1.965 ;
        RECT  0.070 1.355 0.195 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.310 2.505 0.690 ;
        RECT  2.350 1.110 2.505 1.490 ;
        RECT  1.795 0.310 1.850 0.690 ;
        RECT  1.795 1.110 1.850 1.490 ;
        RECT  1.550 0.800 1.800 0.900 ;
        RECT  1.460 0.510 1.550 1.290 ;
        RECT  0.905 0.320 1.520 0.420 ;
        RECT  1.035 0.510 1.460 0.600 ;
        RECT  0.960 1.200 1.460 1.290 ;
        RECT  0.850 1.200 0.960 1.475 ;
        RECT  0.790 0.320 0.905 0.600 ;
        RECT  0.745 0.745 0.810 0.925 ;
        RECT  0.655 0.745 0.745 1.290 ;
        RECT  0.360 1.200 0.655 1.290 ;
        RECT  0.270 0.510 0.360 1.290 ;
        RECT  0.180 0.510 0.270 0.600 ;
        RECT  0.080 0.325 0.180 0.600 ;
    END
END MAOI22D4

MACRO MOAI22D0
    CLASS CORE ;
    FOREIGN MOAI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.290 ;
        RECT  1.040 0.510 1.450 0.600 ;
        RECT  0.965 1.200 1.450 1.290 ;
        RECT  0.850 1.200 0.965 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.565 0.920 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.980 0.710 1.050 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.695 -0.165 1.600 0.165 ;
        RECT  0.575 -0.165 0.695 0.400 ;
        RECT  0.000 -0.165 0.575 0.165 ;
        RECT  0.475 0.290 0.575 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 1.635 1.600 1.965 ;
        RECT  1.395 1.400 1.505 1.965 ;
        RECT  1.295 1.400 1.395 1.510 ;
        RECT  0.705 1.635 1.395 1.965 ;
        RECT  0.595 1.335 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.335 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.905 0.290 1.535 0.400 ;
        RECT  0.790 0.290 0.905 0.480 ;
        RECT  0.745 0.760 0.870 0.870 ;
        RECT  0.655 0.760 0.745 1.245 ;
        RECT  0.445 1.115 0.655 1.245 ;
        RECT  0.360 1.115 0.445 1.490 ;
        RECT  0.335 0.510 0.360 1.490 ;
        RECT  0.270 0.510 0.335 1.245 ;
        RECT  0.185 0.510 0.270 0.600 ;
        RECT  0.075 0.280 0.185 0.600 ;
    END
END MOAI22D0

MACRO MOAI22D1
    CLASS CORE ;
    FOREIGN MOAI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.290 ;
        RECT  1.035 0.510 1.450 0.600 ;
        RECT  0.960 1.200 1.450 1.290 ;
        RECT  0.955 1.200 0.960 1.490 ;
        RECT  0.850 1.045 0.955 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.555 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.090 ;
        RECT  0.970 0.710 1.045 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.680 -0.165 1.600 0.165 ;
        RECT  0.490 -0.165 0.680 0.400 ;
        RECT  0.000 -0.165 0.490 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 1.635 1.600 1.965 ;
        RECT  1.305 1.400 1.485 1.965 ;
        RECT  0.745 1.635 1.305 1.965 ;
        RECT  0.555 1.400 0.745 1.965 ;
        RECT  0.195 1.635 0.555 1.965 ;
        RECT  0.070 1.355 0.195 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.905 0.275 1.490 0.400 ;
        RECT  0.790 0.275 0.905 0.600 ;
        RECT  0.745 0.745 0.810 0.925 ;
        RECT  0.655 0.745 0.745 1.290 ;
        RECT  0.360 1.200 0.655 1.290 ;
        RECT  0.270 0.510 0.360 1.290 ;
        RECT  0.190 0.510 0.270 0.600 ;
        RECT  0.070 0.325 0.190 0.600 ;
    END
END MOAI22D1

MACRO MOAI22D2
    CLASS CORE ;
    FOREIGN MOAI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.955 0.275 2.015 0.675 ;
        RECT  1.955 1.045 2.015 1.490 ;
        RECT  1.900 0.275 1.955 1.490 ;
        RECT  1.845 0.510 1.900 1.195 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.360 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.090 ;
        RECT  0.970 0.710 1.045 0.920 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.565 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 -0.165 2.400 0.165 ;
        RECT  2.160 -0.165 2.275 0.675 ;
        RECT  1.785 -0.165 2.160 0.165 ;
        RECT  1.615 -0.165 1.785 0.405 ;
        RECT  1.485 -0.165 1.615 0.165 ;
        RECT  1.315 -0.165 1.485 0.405 ;
        RECT  0.745 -0.165 1.315 0.165 ;
        RECT  0.555 -0.165 0.745 0.405 ;
        RECT  0.180 -0.165 0.555 0.165 ;
        RECT  0.070 -0.165 0.180 0.530 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 1.635 2.400 1.965 ;
        RECT  2.160 1.045 2.275 1.965 ;
        RECT  1.785 1.635 2.160 1.965 ;
        RECT  1.615 1.395 1.785 1.965 ;
        RECT  0.650 1.635 1.615 1.965 ;
        RECT  0.520 1.240 0.650 1.965 ;
        RECT  0.000 1.635 0.520 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.535 0.510 1.665 1.295 ;
        RECT  0.980 0.510 1.535 0.600 ;
        RECT  1.015 1.205 1.535 1.295 ;
        RECT  0.905 1.395 1.490 1.525 ;
        RECT  0.850 0.360 0.980 0.600 ;
        RECT  0.790 1.205 0.905 1.525 ;
        RECT  0.745 0.750 0.810 0.930 ;
        RECT  0.655 0.510 0.745 0.930 ;
        RECT  0.360 0.510 0.655 0.600 ;
        RECT  0.270 0.510 0.360 1.315 ;
        RECT  0.195 1.200 0.270 1.315 ;
        RECT  0.065 1.200 0.195 1.515 ;
    END
END MOAI22D2

MACRO MOAI22D4
    CLASS CORE ;
    FOREIGN MOAI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.310 2.505 0.690 ;
        RECT  2.250 1.110 2.505 1.490 ;
        RECT  1.950 0.310 2.250 1.490 ;
        RECT  1.845 0.310 1.950 0.690 ;
        RECT  1.845 1.110 1.950 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.555 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.510 1.155 0.890 ;
        RECT  0.950 0.780 1.045 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.565 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.735 -0.165 2.800 0.165 ;
        RECT  2.615 -0.165 2.735 0.690 ;
        RECT  1.655 -0.165 2.615 0.165 ;
        RECT  1.465 -0.165 1.655 0.405 ;
        RECT  0.745 -0.165 1.465 0.165 ;
        RECT  0.555 -0.165 0.745 0.405 ;
        RECT  0.180 -0.165 0.555 0.165 ;
        RECT  0.070 -0.165 0.180 0.600 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.735 1.635 2.800 1.965 ;
        RECT  2.615 1.110 2.735 1.965 ;
        RECT  1.715 1.635 2.615 1.965 ;
        RECT  1.545 1.385 1.715 1.965 ;
        RECT  0.650 1.635 1.545 1.965 ;
        RECT  0.520 1.240 0.650 1.965 ;
        RECT  0.000 1.635 0.520 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.310 2.505 0.690 ;
        RECT  2.350 1.110 2.505 1.490 ;
        RECT  1.650 0.510 1.750 1.295 ;
        RECT  1.355 0.510 1.650 0.600 ;
        RECT  1.200 1.205 1.650 1.295 ;
        RECT  0.920 1.025 1.505 1.115 ;
        RECT  1.265 0.275 1.355 0.600 ;
        RECT  0.955 0.275 1.265 0.365 ;
        RECT  1.070 1.205 1.200 1.515 ;
        RECT  0.850 0.275 0.955 0.600 ;
        RECT  0.790 1.025 0.920 1.515 ;
        RECT  0.745 0.780 0.850 0.890 ;
        RECT  0.655 0.510 0.745 0.890 ;
        RECT  0.360 0.510 0.655 0.600 ;
        RECT  0.270 0.510 0.360 1.315 ;
        RECT  0.190 1.200 0.270 1.315 ;
        RECT  0.065 1.200 0.190 1.515 ;
    END
END MOAI22D4

MACRO MUX2D0
    CLASS CORE ;
    FOREIGN MUX2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.275 1.750 1.315 ;
        RECT  1.615 0.275 1.650 0.485 ;
        RECT  1.615 1.105 1.650 1.315 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.365 1.090 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.710 0.610 0.960 ;
        RECT  0.450 0.710 0.550 1.090 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.400 -0.165 1.800 0.165 ;
        RECT  0.400 0.490 0.500 0.600 ;
        RECT  0.290 -0.165 0.400 0.600 ;
        RECT  0.000 -0.165 0.290 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.505 1.635 1.800 1.965 ;
        RECT  0.335 1.400 0.505 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.505 1.445 1.680 1.545 ;
        RECT  1.395 1.205 1.505 1.545 ;
        RECT  1.010 1.205 1.395 1.295 ;
        RECT  0.955 1.435 1.165 1.545 ;
        RECT  0.890 0.275 1.010 1.295 ;
        RECT  0.710 1.435 0.955 1.525 ;
        RECT  0.620 1.200 0.710 1.525 ;
        RECT  0.175 1.200 0.620 1.290 ;
        RECT  0.155 0.435 0.180 0.625 ;
        RECT  0.155 1.200 0.175 1.505 ;
        RECT  0.065 0.435 0.155 1.505 ;
    END
END MUX2D0

MACRO MUX2D1
    CLASS CORE ;
    FOREIGN MUX2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.835 0.510 1.950 1.525 ;
        RECT  1.825 0.275 1.835 1.525 ;
        RECT  1.730 0.275 1.825 0.650 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.490 1.555 0.900 ;
        RECT  1.350 0.710 1.445 0.900 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0331 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.695 0.600 0.940 ;
        RECT  0.450 0.695 0.550 1.130 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.590 -0.165 2.000 0.165 ;
        RECT  1.400 -0.165 1.590 0.400 ;
        RECT  0.480 -0.165 1.400 0.165 ;
        RECT  0.310 -0.165 0.480 0.575 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.685 1.635 2.000 1.965 ;
        RECT  1.515 1.415 1.685 1.965 ;
        RECT  0.505 1.635 1.515 1.965 ;
        RECT  0.335 1.445 0.505 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.760 1.735 1.325 ;
        RECT  1.170 1.235 1.645 1.325 ;
        RECT  1.250 1.025 1.410 1.145 ;
        RECT  0.765 1.425 1.280 1.525 ;
        RECT  1.150 0.275 1.250 1.145 ;
        RECT  1.010 1.235 1.170 1.335 ;
        RECT  0.960 0.825 1.010 1.335 ;
        RECT  0.920 0.435 0.960 1.335 ;
        RECT  0.870 0.435 0.920 0.915 ;
        RECT  0.780 1.050 0.820 1.155 ;
        RECT  0.690 0.465 0.780 1.155 ;
        RECT  0.675 1.265 0.765 1.525 ;
        RECT  0.570 0.465 0.690 0.575 ;
        RECT  0.640 1.050 0.690 1.155 ;
        RECT  0.175 1.265 0.675 1.355 ;
        RECT  0.160 0.445 0.175 0.615 ;
        RECT  0.160 1.265 0.175 1.515 ;
        RECT  0.065 0.445 0.160 1.515 ;
    END
END MUX2D1

MACRO MUX2D2
    CLASS CORE ;
    FOREIGN MUX2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.510 1.955 1.490 ;
        RECT  1.830 0.510 1.845 0.650 ;
        RECT  1.725 1.300 1.845 1.490 ;
        RECT  1.730 0.275 1.830 0.650 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0679 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.130 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.490 1.555 0.930 ;
        RECT  1.350 0.725 1.445 0.930 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.695 0.600 0.940 ;
        RECT  0.445 0.695 0.550 1.130 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.135 -0.165 2.200 0.165 ;
        RECT  1.945 -0.165 2.135 0.400 ;
        RECT  1.600 -0.165 1.945 0.165 ;
        RECT  1.410 -0.165 1.600 0.400 ;
        RECT  0.480 -0.165 1.410 0.165 ;
        RECT  0.310 -0.165 0.480 0.575 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.505 1.635 2.200 1.965 ;
        RECT  0.335 1.445 0.505 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.760 1.735 1.155 ;
        RECT  1.600 1.055 1.645 1.155 ;
        RECT  1.510 1.055 1.600 1.335 ;
        RECT  1.055 1.245 1.510 1.335 ;
        RECT  1.250 1.055 1.380 1.155 ;
        RECT  1.160 0.275 1.250 1.155 ;
        RECT  0.765 1.425 1.250 1.525 ;
        RECT  0.965 0.825 1.055 1.335 ;
        RECT  0.960 0.825 0.965 0.915 ;
        RECT  0.870 0.435 0.960 0.915 ;
        RECT  0.780 1.050 0.820 1.155 ;
        RECT  0.690 0.465 0.780 1.155 ;
        RECT  0.675 1.265 0.765 1.525 ;
        RECT  0.570 0.465 0.690 0.575 ;
        RECT  0.640 1.050 0.690 1.155 ;
        RECT  0.175 1.265 0.675 1.355 ;
        RECT  0.155 0.445 0.175 0.615 ;
        RECT  0.155 1.265 0.175 1.515 ;
        RECT  0.065 0.445 0.155 1.515 ;
    END
END MUX2D2

MACRO MUX2D4
    CLASS CORE ;
    FOREIGN MUX2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.105 0.690 ;
        RECT  3.050 1.110 3.105 1.490 ;
        RECT  2.750 0.310 3.050 1.490 ;
        RECT  2.450 0.310 2.750 0.690 ;
        RECT  2.450 1.110 2.750 1.490 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0673 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.710 1.755 1.195 ;
        RECT  1.610 0.710 1.645 0.930 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.710 2.155 1.195 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.555 0.890 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.335 -0.165 3.400 0.165 ;
        RECT  3.215 -0.165 3.335 0.690 ;
        RECT  0.480 -0.165 3.215 0.165 ;
        RECT  0.310 -0.165 0.480 0.410 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.335 1.635 3.400 1.965 ;
        RECT  3.215 1.110 3.335 1.965 ;
        RECT  1.800 1.635 3.215 1.965 ;
        RECT  1.610 1.515 1.800 1.965 ;
        RECT  0.480 1.635 1.610 1.965 ;
        RECT  0.310 1.375 0.480 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.450 0.310 2.650 0.690 ;
        RECT  2.450 1.110 2.650 1.490 ;
        RECT  2.340 0.800 2.560 0.910 ;
        RECT  2.245 0.275 2.340 0.910 ;
        RECT  1.000 0.275 2.245 0.365 ;
        RECT  1.935 0.490 2.115 0.600 ;
        RECT  1.935 1.335 2.115 1.425 ;
        RECT  1.845 0.490 1.935 1.425 ;
        RECT  1.250 1.335 1.845 1.425 ;
        RECT  1.400 0.475 1.520 1.195 ;
        RECT  1.340 0.740 1.400 0.930 ;
        RECT  1.150 0.455 1.250 1.425 ;
        RECT  0.865 0.275 1.000 1.320 ;
        RECT  0.595 0.285 0.725 0.600 ;
        RECT  0.595 1.055 0.725 1.525 ;
        RECT  0.200 0.510 0.595 0.600 ;
        RECT  0.200 1.055 0.595 1.145 ;
        RECT  0.150 0.285 0.200 0.600 ;
        RECT  0.150 1.055 0.200 1.525 ;
        RECT  0.060 0.285 0.150 1.525 ;
    END
END MUX2D4

MACRO MUX2ND0
    CLASS CORE ;
    FOREIGN MUX2ND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.215 1.045 1.325 ;
        RECT  0.850 0.435 0.950 1.325 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0667 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.360 1.090 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.510 1.550 0.900 ;
        RECT  1.350 0.710 1.445 0.900 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0328 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.710 0.600 0.940 ;
        RECT  0.450 0.710 0.550 1.090 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.165 1.600 0.165 ;
        RECT  1.270 0.290 1.545 0.400 ;
        RECT  1.140 -0.165 1.270 0.400 ;
        RECT  0.400 -0.165 1.140 0.165 ;
        RECT  0.400 0.490 0.500 0.600 ;
        RECT  0.290 -0.165 0.400 0.600 ;
        RECT  0.000 -0.165 0.290 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 1.635 1.600 1.965 ;
        RECT  1.395 1.040 1.525 1.965 ;
        RECT  0.480 1.635 1.395 1.965 ;
        RECT  0.310 1.380 0.480 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.145 0.775 1.240 1.525 ;
        RECT  1.040 0.775 1.145 0.945 ;
        RECT  0.710 1.435 1.145 1.525 ;
        RECT  0.620 1.200 0.710 1.525 ;
        RECT  0.185 1.200 0.620 1.290 ;
        RECT  0.155 0.445 0.185 0.615 ;
        RECT  0.155 1.200 0.185 1.505 ;
        RECT  0.065 0.445 0.155 1.505 ;
    END
END MUX2ND0

MACRO MUX2ND1
    CLASS CORE ;
    FOREIGN MUX2ND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.275 2.350 1.490 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0679 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.130 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.490 1.555 0.930 ;
        RECT  1.350 0.725 1.445 0.930 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0348 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.695 0.600 0.895 ;
        RECT  0.445 0.695 0.555 1.130 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.590 -0.165 2.400 0.165 ;
        RECT  1.400 -0.165 1.590 0.400 ;
        RECT  0.480 -0.165 1.400 0.165 ;
        RECT  0.310 -0.165 0.480 0.575 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.505 1.635 2.400 1.965 ;
        RECT  0.335 1.445 0.505 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.965 0.510 2.110 1.470 ;
        RECT  1.845 0.510 1.965 0.650 ;
        RECT  1.700 1.305 1.965 1.470 ;
        RECT  1.715 0.265 1.845 0.650 ;
        RECT  1.645 0.760 1.755 1.155 ;
        RECT  1.575 1.055 1.645 1.155 ;
        RECT  1.485 1.055 1.575 1.335 ;
        RECT  1.055 1.245 1.485 1.335 ;
        RECT  1.250 1.055 1.360 1.155 ;
        RECT  0.765 1.425 1.255 1.525 ;
        RECT  1.160 0.275 1.250 1.155 ;
        RECT  0.990 0.805 1.055 1.335 ;
        RECT  0.940 0.435 0.990 1.335 ;
        RECT  0.870 0.435 0.940 0.915 ;
        RECT  0.690 0.465 0.780 1.165 ;
        RECT  0.675 1.265 0.765 1.525 ;
        RECT  0.570 0.465 0.690 0.575 ;
        RECT  0.665 0.985 0.690 1.165 ;
        RECT  0.175 1.265 0.675 1.355 ;
        RECT  0.155 0.445 0.175 0.615 ;
        RECT  0.155 1.265 0.175 1.515 ;
        RECT  0.065 0.445 0.155 1.515 ;
    END
END MUX2ND1

MACRO MUX2ND2
    CLASS CORE ;
    FOREIGN MUX2ND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.275 2.350 1.490 ;
        RECT  2.165 0.275 2.250 0.675 ;
        RECT  2.165 1.045 2.250 1.490 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0565 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.130 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.490 1.555 0.930 ;
        RECT  1.335 0.725 1.445 0.930 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.695 0.585 0.915 ;
        RECT  0.445 0.695 0.555 1.130 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.570 -0.165 2.600 0.165 ;
        RECT  1.380 -0.165 1.570 0.400 ;
        RECT  0.475 -0.165 1.380 0.165 ;
        RECT  0.305 -0.165 0.475 0.575 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 1.635 2.600 1.965 ;
        RECT  0.330 1.445 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.510 2.055 1.465 ;
        RECT  1.810 0.510 1.925 0.650 ;
        RECT  1.650 1.325 1.925 1.465 ;
        RECT  1.685 0.255 1.810 0.650 ;
        RECT  1.645 0.760 1.745 1.155 ;
        RECT  1.555 1.055 1.645 1.155 ;
        RECT  1.465 1.055 1.555 1.335 ;
        RECT  1.030 1.245 1.465 1.335 ;
        RECT  1.245 1.055 1.345 1.155 ;
        RECT  1.140 0.275 1.245 1.155 ;
        RECT  0.760 1.425 1.195 1.525 ;
        RECT  0.980 0.810 1.030 1.335 ;
        RECT  0.920 0.415 0.980 1.335 ;
        RECT  0.865 0.415 0.920 0.915 ;
        RECT  0.685 0.465 0.775 1.175 ;
        RECT  0.670 1.265 0.760 1.525 ;
        RECT  0.565 0.465 0.685 0.575 ;
        RECT  0.650 1.005 0.685 1.175 ;
        RECT  0.180 1.265 0.670 1.355 ;
        RECT  0.155 1.265 0.180 1.515 ;
        RECT  0.155 0.445 0.175 0.615 ;
        RECT  0.065 0.445 0.155 1.515 ;
    END
END MUX2ND2

MACRO MUX2ND4
    CLASS CORE ;
    FOREIGN MUX2ND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.310 3.705 0.690 ;
        RECT  3.650 1.110 3.705 1.490 ;
        RECT  3.350 0.310 3.650 1.490 ;
        RECT  3.020 0.310 3.350 0.690 ;
        RECT  3.020 1.110 3.350 1.490 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0673 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.710 1.755 1.100 ;
        RECT  1.610 0.710 1.645 0.930 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.710 2.155 1.100 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.555 0.890 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.925 -0.165 4.000 0.165 ;
        RECT  3.815 -0.165 3.925 0.690 ;
        RECT  2.890 -0.165 3.815 0.165 ;
        RECT  2.740 -0.165 2.890 0.510 ;
        RECT  0.480 -0.165 2.740 0.165 ;
        RECT  0.310 -0.165 0.480 0.410 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.925 1.635 4.000 1.965 ;
        RECT  3.815 1.110 3.925 1.965 ;
        RECT  2.880 1.635 3.815 1.965 ;
        RECT  2.750 1.295 2.880 1.965 ;
        RECT  2.350 1.635 2.750 1.965 ;
        RECT  2.205 1.295 2.350 1.965 ;
        RECT  1.800 1.635 2.205 1.965 ;
        RECT  1.610 1.515 1.800 1.965 ;
        RECT  0.480 1.635 1.610 1.965 ;
        RECT  0.310 1.375 0.480 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 0.310 3.250 0.690 ;
        RECT  3.020 1.110 3.250 1.490 ;
        RECT  2.810 0.795 3.200 0.905 ;
        RECT  2.700 0.600 2.810 1.205 ;
        RECT  2.605 0.600 2.700 0.710 ;
        RECT  2.605 1.095 2.700 1.205 ;
        RECT  2.495 0.310 2.605 0.710 ;
        RECT  2.495 1.095 2.605 1.505 ;
        RECT  2.360 0.800 2.590 0.900 ;
        RECT  2.265 0.275 2.360 0.900 ;
        RECT  1.000 0.275 2.265 0.365 ;
        RECT  1.935 0.490 2.115 0.600 ;
        RECT  1.935 1.315 2.115 1.425 ;
        RECT  1.845 0.490 1.935 1.425 ;
        RECT  1.250 1.335 1.845 1.425 ;
        RECT  1.420 0.495 1.520 1.195 ;
        RECT  1.340 0.740 1.420 0.930 ;
        RECT  1.150 0.455 1.250 1.425 ;
        RECT  0.865 0.275 1.000 1.320 ;
        RECT  0.595 0.285 0.725 0.600 ;
        RECT  0.595 1.055 0.725 1.525 ;
        RECT  0.200 0.510 0.595 0.600 ;
        RECT  0.200 1.055 0.595 1.145 ;
        RECT  0.150 0.285 0.200 0.600 ;
        RECT  0.150 1.055 0.200 1.525 ;
        RECT  0.060 0.285 0.150 1.525 ;
    END
END MUX2ND4

MACRO MUX3D0
    CLASS CORE ;
    FOREIGN MUX3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.435 3.150 1.490 ;
        RECT  3.025 0.435 3.050 0.645 ;
        RECT  3.015 1.265 3.050 1.490 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.710 1.750 1.090 ;
        RECT  1.605 0.710 1.640 0.930 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0559 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.355 1.090 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 0.710 2.755 1.090 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.110 1.550 1.490 ;
        RECT  1.425 0.780 1.515 1.490 ;
        RECT  1.300 0.780 1.425 0.890 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.710 0.585 0.915 ;
        RECT  0.450 0.710 0.550 1.090 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.480 -0.165 3.200 0.165 ;
        RECT  0.310 -0.165 0.480 0.595 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.865 1.635 3.200 1.965 ;
        RECT  2.755 1.280 2.865 1.965 ;
        RECT  0.500 1.635 2.755 1.965 ;
        RECT  0.330 1.445 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.935 0.835 2.960 1.035 ;
        RECT  2.845 0.290 2.935 1.035 ;
        RECT  2.335 0.290 2.845 0.380 ;
        RECT  2.525 1.330 2.655 1.440 ;
        RECT  2.525 0.490 2.625 0.600 ;
        RECT  2.425 0.490 2.525 1.440 ;
        RECT  2.215 0.290 2.335 1.490 ;
        RECT  2.035 0.275 2.125 1.490 ;
        RECT  0.965 0.275 2.035 0.375 ;
        RECT  1.935 1.375 2.035 1.490 ;
        RECT  1.855 0.520 1.945 1.285 ;
        RECT  1.640 0.520 1.855 0.620 ;
        RECT  1.670 1.180 1.855 1.285 ;
        RECT  1.210 0.520 1.350 0.630 ;
        RECT  1.210 1.165 1.335 1.275 ;
        RECT  0.760 1.425 1.235 1.525 ;
        RECT  1.120 0.520 1.210 1.275 ;
        RECT  0.965 0.825 1.030 1.315 ;
        RECT  0.930 0.275 0.965 1.315 ;
        RECT  0.865 0.275 0.930 0.915 ;
        RECT  0.685 0.485 0.775 1.175 ;
        RECT  0.670 1.265 0.760 1.525 ;
        RECT  0.570 0.485 0.685 0.595 ;
        RECT  0.650 1.005 0.685 1.175 ;
        RECT  0.180 1.265 0.670 1.355 ;
        RECT  0.140 0.495 0.220 0.605 ;
        RECT  0.140 1.265 0.180 1.515 ;
        RECT  0.050 0.495 0.140 1.515 ;
    END
END MUX3D0

MACRO MUX3D1
    CLASS CORE ;
    FOREIGN MUX3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.310 3.150 1.490 ;
        RECT  3.025 0.310 3.050 0.600 ;
        RECT  3.025 1.045 3.050 1.490 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0636 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.710 1.755 1.090 ;
        RECT  1.605 0.710 1.640 0.930 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0679 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.130 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.645 0.710 2.755 1.290 ;
        RECT  2.620 0.710 2.645 0.930 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.110 1.550 1.490 ;
        RECT  1.425 0.755 1.515 1.490 ;
        RECT  1.300 0.755 1.425 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.695 0.585 0.915 ;
        RECT  0.450 0.695 0.550 1.130 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.475 -0.165 3.200 0.165 ;
        RECT  0.305 -0.165 0.475 0.575 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.635 3.200 1.965 ;
        RECT  2.725 1.380 2.900 1.965 ;
        RECT  0.500 1.635 2.725 1.965 ;
        RECT  0.330 1.445 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.935 0.740 2.960 0.930 ;
        RECT  2.845 0.275 2.935 0.930 ;
        RECT  2.335 0.275 2.845 0.365 ;
        RECT  2.525 1.380 2.635 1.490 ;
        RECT  2.525 0.475 2.625 0.600 ;
        RECT  2.425 0.475 2.525 1.490 ;
        RECT  2.215 0.275 2.335 1.490 ;
        RECT  2.035 0.275 2.125 1.490 ;
        RECT  0.970 0.275 2.035 0.385 ;
        RECT  1.935 1.380 2.035 1.490 ;
        RECT  1.855 0.510 1.945 1.290 ;
        RECT  1.640 0.510 1.855 0.620 ;
        RECT  1.690 1.180 1.855 1.290 ;
        RECT  1.210 0.495 1.345 0.605 ;
        RECT  1.210 1.100 1.335 1.270 ;
        RECT  0.760 1.425 1.235 1.525 ;
        RECT  1.120 0.495 1.210 1.270 ;
        RECT  0.970 0.825 1.030 1.315 ;
        RECT  0.920 0.275 0.970 1.315 ;
        RECT  0.865 0.275 0.920 0.915 ;
        RECT  0.685 0.465 0.775 1.175 ;
        RECT  0.670 1.265 0.760 1.525 ;
        RECT  0.565 0.465 0.685 0.575 ;
        RECT  0.650 1.005 0.685 1.175 ;
        RECT  0.180 1.265 0.670 1.355 ;
        RECT  0.155 1.265 0.180 1.515 ;
        RECT  0.155 0.445 0.175 0.615 ;
        RECT  0.065 0.445 0.155 1.515 ;
    END
END MUX3D1

MACRO MUX3D2
    CLASS CORE ;
    FOREIGN MUX3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.295 3.150 1.490 ;
        RECT  2.935 0.295 3.050 0.420 ;
        RECT  2.965 1.045 3.050 1.490 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0636 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.710 1.755 1.090 ;
        RECT  1.605 0.710 1.640 0.930 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0565 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.130 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.645 0.710 2.760 1.290 ;
        RECT  2.620 0.710 2.645 0.930 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 1.110 1.550 1.490 ;
        RECT  1.425 0.785 1.515 1.490 ;
        RECT  1.300 0.785 1.425 0.885 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.695 0.585 0.915 ;
        RECT  0.450 0.695 0.550 1.130 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.475 -0.165 3.400 0.165 ;
        RECT  0.305 -0.165 0.475 0.575 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 1.635 3.400 1.965 ;
        RECT  0.330 1.445 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.870 0.510 2.960 0.930 ;
        RECT  2.825 0.510 2.870 0.600 ;
        RECT  2.735 0.275 2.825 0.600 ;
        RECT  2.315 0.275 2.735 0.365 ;
        RECT  2.525 0.505 2.625 0.620 ;
        RECT  2.525 1.380 2.615 1.490 ;
        RECT  2.425 0.505 2.525 1.490 ;
        RECT  2.215 0.275 2.315 1.490 ;
        RECT  2.035 0.275 2.125 1.490 ;
        RECT  0.985 0.275 2.035 0.385 ;
        RECT  1.905 1.380 2.035 1.490 ;
        RECT  1.855 0.510 1.945 1.290 ;
        RECT  1.640 0.510 1.855 0.620 ;
        RECT  1.660 1.180 1.855 1.290 ;
        RECT  1.210 0.505 1.345 0.620 ;
        RECT  1.210 1.170 1.335 1.270 ;
        RECT  1.120 0.505 1.210 1.270 ;
        RECT  0.760 1.425 1.185 1.525 ;
        RECT  0.985 0.805 1.030 1.315 ;
        RECT  0.915 0.275 0.985 1.315 ;
        RECT  0.865 0.275 0.915 0.915 ;
        RECT  0.685 0.465 0.775 1.175 ;
        RECT  0.670 1.265 0.760 1.525 ;
        RECT  0.565 0.465 0.685 0.575 ;
        RECT  0.650 1.005 0.685 1.175 ;
        RECT  0.180 1.265 0.670 1.355 ;
        RECT  0.155 1.265 0.180 1.515 ;
        RECT  0.155 0.445 0.175 0.615 ;
        RECT  0.065 0.445 0.155 1.515 ;
    END
END MUX3D2

MACRO MUX3D4
    CLASS CORE ;
    FOREIGN MUX3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.310 4.905 0.690 ;
        RECT  4.850 1.110 4.905 1.490 ;
        RECT  4.550 0.310 4.850 1.490 ;
        RECT  4.250 0.310 4.550 0.690 ;
        RECT  4.250 1.110 4.550 1.490 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.445 0.710 3.555 1.195 ;
        RECT  3.410 0.710 3.445 0.930 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0679 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.710 1.755 1.195 ;
        RECT  1.595 0.710 1.645 0.930 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.845 0.710 3.955 1.195 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.710 2.155 1.195 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.555 0.890 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.135 -0.165 5.200 0.165 ;
        RECT  5.015 -0.165 5.135 0.690 ;
        RECT  0.475 -0.165 5.015 0.165 ;
        RECT  0.305 -0.165 0.475 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.135 1.635 5.200 1.965 ;
        RECT  5.015 1.110 5.135 1.965 ;
        RECT  3.600 1.635 5.015 1.965 ;
        RECT  3.410 1.505 3.600 1.965 ;
        RECT  1.775 1.635 3.410 1.965 ;
        RECT  1.580 1.505 1.775 1.965 ;
        RECT  0.475 1.635 1.580 1.965 ;
        RECT  0.305 1.375 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.250 0.310 4.450 0.690 ;
        RECT  4.250 1.110 4.450 1.490 ;
        RECT  4.140 0.800 4.360 0.900 ;
        RECT  4.045 0.275 4.140 0.900 ;
        RECT  2.790 0.275 4.045 0.365 ;
        RECT  3.735 0.485 3.915 0.600 ;
        RECT  3.735 1.325 3.915 1.415 ;
        RECT  3.645 0.485 3.735 1.415 ;
        RECT  3.050 1.325 3.645 1.415 ;
        RECT  3.205 0.495 3.320 1.195 ;
        RECT  3.200 0.740 3.205 1.195 ;
        RECT  3.140 0.740 3.200 0.930 ;
        RECT  2.930 0.455 3.050 1.415 ;
        RECT  2.660 0.275 2.790 1.340 ;
        RECT  2.405 0.275 2.535 1.515 ;
        RECT  0.980 0.275 2.405 0.365 ;
        RECT  1.935 0.490 2.090 0.600 ;
        RECT  1.935 1.325 2.085 1.415 ;
        RECT  1.845 0.490 1.935 1.415 ;
        RECT  1.240 1.325 1.845 1.415 ;
        RECT  1.395 0.475 1.505 1.195 ;
        RECT  1.390 0.740 1.395 1.195 ;
        RECT  1.330 0.740 1.390 0.930 ;
        RECT  1.120 0.455 1.240 1.415 ;
        RECT  0.850 0.275 0.980 1.320 ;
        RECT  0.585 0.285 0.715 0.600 ;
        RECT  0.585 1.055 0.715 1.525 ;
        RECT  0.195 0.510 0.585 0.600 ;
        RECT  0.195 1.055 0.585 1.145 ;
        RECT  0.155 0.285 0.195 0.600 ;
        RECT  0.155 1.055 0.195 1.525 ;
        RECT  0.065 0.285 0.155 1.525 ;
    END
END MUX3D4

MACRO MUX3ND0
    CLASS CORE ;
    FOREIGN MUX3ND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0980 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.550 1.210 ;
        RECT  2.405 0.710 2.450 0.800 ;
        RECT  2.405 1.100 2.450 1.210 ;
        RECT  2.295 0.480 2.405 0.800 ;
        RECT  2.295 1.100 2.405 1.465 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0689 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.710 1.765 1.090 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.360 1.110 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0558 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.820 0.710 2.950 1.090 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.510 1.550 0.900 ;
        RECT  1.350 0.710 1.445 0.900 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0331 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.710 0.600 0.960 ;
        RECT  0.450 0.710 0.550 1.090 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.925 -0.165 3.000 0.165 ;
        RECT  2.820 -0.165 2.925 0.585 ;
        RECT  1.595 -0.165 2.820 0.165 ;
        RECT  1.385 -0.165 1.595 0.400 ;
        RECT  0.480 -0.165 1.385 0.165 ;
        RECT  0.370 -0.165 0.480 0.600 ;
        RECT  0.000 -0.165 0.370 0.165 ;
        RECT  0.290 0.490 0.370 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.925 1.635 3.000 1.965 ;
        RECT  2.820 1.200 2.925 1.965 ;
        RECT  1.725 1.635 2.820 1.965 ;
        RECT  1.555 1.490 1.725 1.965 ;
        RECT  0.505 1.635 1.555 1.965 ;
        RECT  0.335 1.445 0.505 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.640 0.490 2.730 1.430 ;
        RECT  2.520 0.490 2.640 0.600 ;
        RECT  2.505 1.320 2.640 1.430 ;
        RECT  2.115 0.255 2.205 1.520 ;
        RECT  1.945 0.255 2.115 0.370 ;
        RECT  2.005 1.290 2.115 1.520 ;
        RECT  1.895 0.480 2.025 1.155 ;
        RECT  1.520 1.290 2.005 1.380 ;
        RECT  1.675 0.480 1.895 0.590 ;
        RECT  1.430 1.205 1.520 1.380 ;
        RECT  0.990 1.205 1.430 1.295 ;
        RECT  1.250 1.015 1.405 1.115 ;
        RECT  1.090 1.405 1.280 1.545 ;
        RECT  1.135 0.265 1.250 1.115 ;
        RECT  0.765 1.405 1.090 1.495 ;
        RECT  0.900 0.435 0.990 1.295 ;
        RECT  0.870 0.435 0.900 0.645 ;
        RECT  0.780 1.055 0.810 1.155 ;
        RECT  0.690 0.465 0.780 1.155 ;
        RECT  0.675 1.265 0.765 1.495 ;
        RECT  0.570 0.465 0.690 0.575 ;
        RECT  0.640 1.055 0.690 1.155 ;
        RECT  0.185 1.265 0.675 1.355 ;
        RECT  0.160 1.265 0.185 1.505 ;
        RECT  0.160 0.425 0.180 0.615 ;
        RECT  0.065 0.425 0.160 1.505 ;
    END
END MUX3ND0

MACRO MUX3ND1
    CLASS CORE ;
    FOREIGN MUX3ND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.420 0.275 3.550 1.490 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0624 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.710 1.750 1.090 ;
        RECT  1.590 0.800 1.640 0.990 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0562 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.125 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.645 0.710 2.755 1.290 ;
        RECT  2.605 0.710 2.645 0.930 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.500 0.510 1.550 0.690 ;
        RECT  1.500 1.110 1.550 1.290 ;
        RECT  1.410 0.510 1.500 1.290 ;
        RECT  1.285 0.780 1.410 0.895 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0349 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.695 0.585 0.885 ;
        RECT  0.450 0.695 0.550 1.125 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.475 -0.165 3.600 0.165 ;
        RECT  0.305 -0.165 0.475 0.575 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 1.635 3.600 1.965 ;
        RECT  0.295 1.415 0.485 1.965 ;
        RECT  0.000 1.635 0.295 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.165 0.305 3.310 1.205 ;
        RECT  2.905 0.305 3.165 0.420 ;
        RECT  3.070 1.045 3.165 1.205 ;
        RECT  2.920 1.045 3.070 1.490 ;
        RECT  2.865 0.510 2.970 0.940 ;
        RECT  2.795 0.510 2.865 0.600 ;
        RECT  2.705 0.275 2.795 0.600 ;
        RECT  2.290 0.275 2.705 0.365 ;
        RECT  2.500 1.380 2.600 1.510 ;
        RECT  2.500 0.495 2.595 0.620 ;
        RECT  2.400 0.495 2.500 1.510 ;
        RECT  2.180 0.275 2.290 1.490 ;
        RECT  1.320 1.380 2.080 1.490 ;
        RECT  0.955 0.275 2.055 0.365 ;
        RECT  1.840 0.510 1.930 1.290 ;
        RECT  1.640 0.510 1.840 0.620 ;
        RECT  1.640 1.180 1.840 1.290 ;
        RECT  1.195 1.005 1.320 1.115 ;
        RECT  1.230 1.205 1.320 1.490 ;
        RECT  1.195 0.510 1.300 0.690 ;
        RECT  0.955 1.205 1.230 1.305 ;
        RECT  1.105 0.510 1.195 1.115 ;
        RECT  0.775 1.415 1.140 1.525 ;
        RECT  0.865 0.275 0.955 1.305 ;
        RECT  0.685 0.465 0.775 1.145 ;
        RECT  0.685 1.235 0.775 1.525 ;
        RECT  0.565 0.465 0.685 0.575 ;
        RECT  0.640 0.975 0.685 1.145 ;
        RECT  0.185 1.235 0.685 1.325 ;
        RECT  0.155 0.445 0.185 0.615 ;
        RECT  0.155 1.235 0.185 1.525 ;
        RECT  0.065 0.445 0.155 1.525 ;
    END
END MUX3ND1

MACRO MUX3ND2
    CLASS CORE ;
    FOREIGN MUX3ND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.545 3.750 1.195 ;
        RECT  3.650 0.275 3.675 1.490 ;
        RECT  3.545 0.275 3.650 0.675 ;
        RECT  3.545 1.045 3.650 1.490 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0635 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.755 1.755 1.290 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.355 1.115 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.750 2.955 1.290 ;
        RECT  2.720 0.750 2.845 0.920 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0557 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.755 1.550 1.290 ;
        RECT  1.400 0.755 1.445 0.945 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0346 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.710 0.620 0.915 ;
        RECT  0.445 0.710 0.555 1.115 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.930 -0.165 4.000 0.165 ;
        RECT  3.810 -0.165 3.930 0.455 ;
        RECT  1.645 -0.165 3.810 0.165 ;
        RECT  1.475 -0.165 1.645 0.285 ;
        RECT  0.475 -0.165 1.475 0.165 ;
        RECT  0.305 -0.165 0.475 0.585 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.635 4.000 1.965 ;
        RECT  3.810 1.330 3.930 1.965 ;
        RECT  1.665 1.635 3.810 1.965 ;
        RECT  1.495 1.405 1.665 1.965 ;
        RECT  0.475 1.635 1.495 1.965 ;
        RECT  0.305 1.410 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.310 0.330 3.430 1.185 ;
        RECT  3.020 0.330 3.310 0.440 ;
        RECT  3.185 1.045 3.310 1.185 ;
        RECT  3.065 1.045 3.185 1.490 ;
        RECT  3.045 0.550 3.135 0.930 ;
        RECT  2.920 0.550 3.045 0.640 ;
        RECT  2.830 0.275 2.920 0.640 ;
        RECT  2.420 0.275 2.830 0.365 ;
        RECT  2.610 0.480 2.720 0.660 ;
        RECT  2.610 1.300 2.720 1.515 ;
        RECT  2.510 0.480 2.610 1.515 ;
        RECT  2.310 0.275 2.420 1.515 ;
        RECT  2.105 0.375 2.200 1.515 ;
        RECT  2.045 0.375 2.105 0.670 ;
        RECT  2.045 1.300 2.105 1.515 ;
        RECT  1.010 0.375 2.045 0.465 ;
        RECT  1.935 0.800 2.015 0.970 ;
        RECT  1.845 0.555 1.935 1.515 ;
        RECT  1.685 0.555 1.845 0.645 ;
        RECT  1.760 1.405 1.845 1.515 ;
        RECT  1.285 0.555 1.380 0.665 ;
        RECT  1.285 1.090 1.335 1.315 ;
        RECT  1.190 0.555 1.285 1.315 ;
        RECT  0.790 1.425 1.270 1.525 ;
        RECT  1.010 1.150 1.080 1.330 ;
        RECT  0.920 0.375 1.010 1.330 ;
        RECT  0.900 0.375 0.920 0.790 ;
        RECT  0.810 0.905 0.825 1.115 ;
        RECT  0.720 0.480 0.810 1.115 ;
        RECT  0.700 1.225 0.790 1.525 ;
        RECT  0.565 0.480 0.720 0.590 ;
        RECT  0.645 1.025 0.720 1.115 ;
        RECT  0.175 1.225 0.700 1.320 ;
        RECT  0.155 0.445 0.175 0.615 ;
        RECT  0.155 1.225 0.175 1.430 ;
        RECT  0.065 0.445 0.155 1.430 ;
    END
END MUX3ND2

MACRO MUX3ND4
    CLASS CORE ;
    FOREIGN MUX3ND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.310 5.305 0.690 ;
        RECT  5.250 1.110 5.305 1.490 ;
        RECT  4.950 0.310 5.250 1.490 ;
        RECT  4.650 0.310 4.950 0.690 ;
        RECT  4.650 1.110 4.950 1.490 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0679 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.820 0.710 3.955 1.195 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0676 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.605 0.710 1.755 1.090 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.710 4.355 1.195 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.710 2.355 0.890 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.1095 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.555 0.890 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.535 -0.165 5.600 0.165 ;
        RECT  5.415 -0.165 5.535 0.690 ;
        RECT  2.355 -0.165 5.415 0.165 ;
        RECT  2.215 -0.165 2.355 0.590 ;
        RECT  0.485 -0.165 2.215 0.165 ;
        RECT  0.315 -0.165 0.485 0.405 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.535 1.635 5.600 1.965 ;
        RECT  5.415 1.110 5.535 1.965 ;
        RECT  4.000 1.635 5.415 1.965 ;
        RECT  3.810 1.515 4.000 1.965 ;
        RECT  1.795 1.635 3.810 1.965 ;
        RECT  1.625 1.505 1.795 1.965 ;
        RECT  0.485 1.635 1.625 1.965 ;
        RECT  0.315 1.290 0.485 1.965 ;
        RECT  0.000 1.635 0.315 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.650 0.310 4.850 0.690 ;
        RECT  4.650 1.110 4.850 1.490 ;
        RECT  4.540 0.800 4.770 0.900 ;
        RECT  4.445 0.275 4.540 0.900 ;
        RECT  2.650 0.275 4.445 0.365 ;
        RECT  4.135 0.490 4.315 0.600 ;
        RECT  4.135 1.335 4.315 1.425 ;
        RECT  4.045 0.490 4.135 1.425 ;
        RECT  3.400 1.335 4.045 1.425 ;
        RECT  3.635 0.495 3.730 1.195 ;
        RECT  3.505 0.745 3.635 0.935 ;
        RECT  3.400 0.455 3.510 0.625 ;
        RECT  3.290 0.455 3.400 1.425 ;
        RECT  3.050 0.495 3.165 1.525 ;
        RECT  2.575 1.435 3.050 1.525 ;
        RECT  2.790 0.495 2.885 1.345 ;
        RECT  2.320 1.255 2.790 1.345 ;
        RECT  2.560 0.275 2.650 1.155 ;
        RECT  2.510 0.275 2.560 0.685 ;
        RECT  2.405 1.045 2.560 1.155 ;
        RECT  2.230 1.255 2.320 1.415 ;
        RECT  0.990 1.325 2.230 1.415 ;
        RECT  1.935 0.435 2.105 0.565 ;
        RECT  1.935 1.095 2.095 1.215 ;
        RECT  1.845 0.325 1.935 1.215 ;
        RECT  1.175 0.325 1.845 0.415 ;
        RECT  1.400 0.505 1.510 1.175 ;
        RECT  1.385 0.505 1.400 0.920 ;
        RECT  1.285 0.750 1.385 0.920 ;
        RECT  1.175 1.085 1.290 1.215 ;
        RECT  1.080 0.325 1.175 1.215 ;
        RECT  0.860 0.285 0.990 1.415 ;
        RECT  0.595 0.285 0.725 0.600 ;
        RECT  0.595 1.055 0.725 1.525 ;
        RECT  0.205 0.510 0.595 0.600 ;
        RECT  0.205 1.055 0.595 1.170 ;
        RECT  0.155 0.285 0.205 0.600 ;
        RECT  0.155 1.055 0.205 1.525 ;
        RECT  0.065 0.285 0.155 1.525 ;
    END
END MUX3ND4

MACRO MUX4D0
    CLASS CORE ;
    FOREIGN MUX4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.310 4.550 1.400 ;
        RECT  4.425 0.310 4.450 0.655 ;
        RECT  4.425 1.100 4.450 1.400 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0527 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.710 4.155 1.090 ;
        RECT  4.020 0.710 4.045 0.930 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0833 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.710 1.750 1.090 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.090 ;
        RECT  1.095 0.710 1.245 0.925 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.705 2.955 1.090 ;
        RECT  2.775 0.705 2.845 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0266 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 1.965 1.090 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.165 4.600 0.165 ;
        RECT  1.655 -0.165 1.765 0.395 ;
        RECT  1.430 -0.165 1.655 0.165 ;
        RECT  1.285 -0.165 1.430 0.395 ;
        RECT  0.195 -0.165 1.285 0.165 ;
        RECT  0.065 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.635 4.600 1.965 ;
        RECT  1.690 1.445 1.860 1.965 ;
        RECT  1.305 1.635 1.690 1.965 ;
        RECT  1.135 1.445 1.305 1.965 ;
        RECT  0.185 1.635 1.135 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.335 0.810 4.360 0.990 ;
        RECT  4.245 0.810 4.335 1.525 ;
        RECT  3.455 1.435 4.245 1.525 ;
        RECT  3.930 0.375 4.055 0.545 ;
        RECT  3.930 1.235 4.045 1.345 ;
        RECT  3.840 0.375 3.930 1.345 ;
        RECT  3.725 0.780 3.840 0.970 ;
        RECT  3.635 1.220 3.730 1.345 ;
        RECT  3.635 0.275 3.715 0.645 ;
        RECT  3.545 0.275 3.635 1.345 ;
        RECT  2.445 0.275 3.545 0.365 ;
        RECT  3.335 0.455 3.455 1.525 ;
        RECT  3.075 0.455 3.200 1.525 ;
        RECT  2.170 1.435 3.075 1.525 ;
        RECT  2.655 0.475 2.770 0.585 ;
        RECT  2.655 1.235 2.755 1.345 ;
        RECT  2.565 0.475 2.655 1.345 ;
        RECT  2.345 0.275 2.445 1.345 ;
        RECT  1.945 0.315 2.255 0.425 ;
        RECT  2.060 1.265 2.170 1.525 ;
        RECT  2.055 0.515 2.165 1.175 ;
        RECT  0.725 1.265 2.060 1.355 ;
        RECT  1.855 0.315 1.945 0.600 ;
        RECT  1.535 0.505 1.855 0.600 ;
        RECT  1.445 0.505 1.535 1.155 ;
        RECT  1.195 0.505 1.445 0.615 ;
        RECT  1.095 0.315 1.195 0.615 ;
        RECT  0.710 0.315 1.095 0.425 ;
        RECT  0.875 0.515 0.985 1.175 ;
        RECT  0.605 0.515 0.725 1.355 ;
        RECT  0.335 0.275 0.445 1.355 ;
    END
END MUX4D0

MACRO MUX4D1
    CLASS CORE ;
    FOREIGN MUX4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.275 4.550 1.525 ;
        RECT  4.425 0.275 4.450 0.675 ;
        RECT  4.425 1.045 4.450 1.525 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0661 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.710 4.155 1.090 ;
        RECT  4.020 0.710 4.045 0.930 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.1045 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.710 1.750 1.090 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0327 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.090 ;
        RECT  1.095 0.710 1.245 0.925 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.705 2.955 1.090 ;
        RECT  2.775 0.705 2.845 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 1.965 1.090 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.165 4.600 0.165 ;
        RECT  1.655 -0.165 1.765 0.395 ;
        RECT  1.430 -0.165 1.655 0.165 ;
        RECT  1.300 -0.165 1.430 0.395 ;
        RECT  0.195 -0.165 1.300 0.165 ;
        RECT  0.065 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.635 4.600 1.965 ;
        RECT  1.690 1.445 1.860 1.965 ;
        RECT  1.305 1.635 1.690 1.965 ;
        RECT  1.135 1.445 1.305 1.965 ;
        RECT  0.195 1.635 1.135 1.965 ;
        RECT  0.065 1.200 0.195 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.335 0.750 4.360 0.930 ;
        RECT  4.245 0.750 4.335 1.525 ;
        RECT  3.455 1.435 4.245 1.525 ;
        RECT  3.930 0.495 4.045 0.600 ;
        RECT  3.930 1.235 4.045 1.345 ;
        RECT  3.840 0.495 3.930 1.345 ;
        RECT  3.725 0.780 3.840 0.970 ;
        RECT  3.635 1.240 3.730 1.345 ;
        RECT  3.635 0.275 3.715 0.645 ;
        RECT  3.545 0.275 3.635 1.345 ;
        RECT  2.445 0.275 3.545 0.365 ;
        RECT  3.335 0.455 3.455 1.525 ;
        RECT  3.075 0.455 3.200 1.525 ;
        RECT  2.170 1.435 3.075 1.525 ;
        RECT  2.655 0.475 2.770 0.585 ;
        RECT  2.655 1.235 2.755 1.345 ;
        RECT  2.565 0.475 2.655 1.345 ;
        RECT  2.345 0.275 2.445 1.345 ;
        RECT  1.945 0.315 2.255 0.425 ;
        RECT  2.060 1.265 2.170 1.525 ;
        RECT  2.055 0.515 2.165 1.175 ;
        RECT  0.725 1.265 2.060 1.355 ;
        RECT  1.855 0.315 1.945 0.600 ;
        RECT  1.535 0.505 1.855 0.600 ;
        RECT  1.445 0.505 1.535 1.155 ;
        RECT  1.195 0.505 1.445 0.615 ;
        RECT  1.095 0.315 1.195 0.615 ;
        RECT  0.705 0.315 1.095 0.425 ;
        RECT  0.875 0.515 0.985 1.175 ;
        RECT  0.605 0.515 0.725 1.355 ;
        RECT  0.335 0.275 0.445 1.355 ;
    END
END MUX4D1

MACRO MUX4D2
    CLASS CORE ;
    FOREIGN MUX4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.275 6.150 1.490 ;
        RECT  5.930 0.275 6.050 0.675 ;
        RECT  5.850 1.110 6.050 1.490 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0669 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.555 0.710 4.630 0.895 ;
        RECT  4.450 0.710 4.555 1.090 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0860 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.435 3.250 1.525 ;
        RECT  1.230 1.255 1.320 1.525 ;
        RECT  0.430 1.255 1.230 1.345 ;
        RECT  0.355 1.020 0.430 1.345 ;
        RECT  0.340 0.700 0.355 1.345 ;
        RECT  0.240 0.700 0.340 1.110 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.710 4.355 0.890 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.710 2.755 0.890 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.755 0.815 0.890 ;
        RECT  0.445 0.510 0.555 0.890 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.710 2.355 0.890 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 6.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 6.400 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.800 0.785 5.940 0.915 ;
        RECT  5.685 0.275 5.800 0.915 ;
        RECT  5.325 0.275 5.685 0.365 ;
        RECT  5.465 0.475 5.595 1.525 ;
        RECT  3.460 1.435 5.465 1.525 ;
        RECT  5.195 0.275 5.325 1.320 ;
        RECT  4.970 0.275 5.075 1.320 ;
        RECT  4.935 0.275 4.970 0.625 ;
        RECT  4.935 1.075 4.970 1.320 ;
        RECT  3.560 0.275 4.935 0.365 ;
        RECT  4.825 0.750 4.880 0.920 ;
        RECT  4.735 0.495 4.825 1.185 ;
        RECT  4.625 0.495 4.735 0.600 ;
        RECT  4.645 1.060 4.735 1.185 ;
        RECT  3.775 1.195 4.355 1.325 ;
        RECT  3.775 0.475 4.345 0.585 ;
        RECT  3.670 0.475 3.775 1.325 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.370 1.255 3.460 1.525 ;
        RECT  3.330 1.075 3.440 1.165 ;
        RECT  1.530 1.255 3.370 1.345 ;
        RECT  2.995 0.475 3.340 0.585 ;
        RECT  3.160 0.255 3.330 0.365 ;
        RECT  2.995 1.055 3.220 1.165 ;
        RECT  1.670 0.275 3.160 0.365 ;
        RECT  2.905 0.475 2.995 1.165 ;
        RECT  2.595 0.475 2.905 0.585 ;
        RECT  2.555 1.055 2.905 1.165 ;
        RECT  1.750 0.475 2.305 0.580 ;
        RECT  1.750 1.055 2.265 1.165 ;
        RECT  1.640 0.475 1.750 1.165 ;
        RECT  1.460 0.255 1.670 0.365 ;
        RECT  1.530 0.475 1.545 0.565 ;
        RECT  1.440 0.475 1.530 1.345 ;
        RECT  0.195 0.275 1.460 0.365 ;
        RECT  1.375 0.475 1.440 0.565 ;
        RECT  1.435 1.075 1.440 1.345 ;
        RECT  1.300 1.075 1.435 1.165 ;
        RECT  1.050 0.475 1.285 0.565 ;
        RECT  1.050 1.075 1.190 1.165 ;
        RECT  0.195 1.435 1.120 1.525 ;
        RECT  0.960 0.475 1.050 1.165 ;
        RECT  0.740 0.475 0.960 0.565 ;
        RECT  0.545 1.075 0.960 1.165 ;
        RECT  0.650 0.475 0.740 0.645 ;
        RECT  0.140 0.275 0.195 0.560 ;
        RECT  0.140 1.220 0.195 1.525 ;
        RECT  0.050 0.275 0.140 1.525 ;
    END
END MUX4D2

MACRO MUX4D4
    CLASS CORE ;
    FOREIGN MUX4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.545 0.275 6.675 0.675 ;
        RECT  6.545 1.035 6.675 1.490 ;
        RECT  6.450 0.520 6.545 0.675 ;
        RECT  6.450 1.035 6.545 1.205 ;
        RECT  6.150 0.520 6.450 1.205 ;
        RECT  6.115 0.520 6.150 0.675 ;
        RECT  6.120 1.035 6.150 1.205 ;
        RECT  5.985 1.035 6.120 1.490 ;
        RECT  5.985 0.275 6.115 0.675 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0669 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.555 0.710 4.630 0.895 ;
        RECT  4.450 0.710 4.555 1.090 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0860 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.435 3.250 1.525 ;
        RECT  1.230 1.255 1.320 1.525 ;
        RECT  0.430 1.255 1.230 1.345 ;
        RECT  0.355 1.020 0.430 1.345 ;
        RECT  0.340 0.700 0.355 1.345 ;
        RECT  0.240 0.700 0.340 1.110 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.710 4.355 0.890 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.710 2.755 0.890 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.755 0.815 0.890 ;
        RECT  0.445 0.510 0.555 0.890 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.710 2.355 0.890 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.935 -0.165 7.000 0.165 ;
        RECT  6.815 -0.165 6.935 0.690 ;
        RECT  6.425 -0.165 6.815 0.165 ;
        RECT  6.235 -0.165 6.425 0.420 ;
        RECT  0.000 -0.165 6.235 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.935 1.635 7.000 1.965 ;
        RECT  6.815 1.110 6.935 1.965 ;
        RECT  6.395 1.635 6.815 1.965 ;
        RECT  6.265 1.325 6.395 1.965 ;
        RECT  5.855 1.635 6.265 1.965 ;
        RECT  5.725 1.085 5.855 1.965 ;
        RECT  0.000 1.635 5.725 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.550 0.275 6.675 0.675 ;
        RECT  6.550 1.035 6.675 1.490 ;
        RECT  5.985 0.275 6.050 0.675 ;
        RECT  5.985 1.035 6.050 1.490 ;
        RECT  5.835 0.785 6.040 0.915 ;
        RECT  5.720 0.275 5.835 0.915 ;
        RECT  5.325 0.275 5.720 0.365 ;
        RECT  5.465 0.475 5.595 1.525 ;
        RECT  3.460 1.435 5.465 1.525 ;
        RECT  5.195 0.275 5.325 1.320 ;
        RECT  4.970 0.275 5.075 1.320 ;
        RECT  4.935 0.275 4.970 0.625 ;
        RECT  4.935 1.075 4.970 1.320 ;
        RECT  3.560 0.275 4.935 0.365 ;
        RECT  4.825 0.750 4.880 0.920 ;
        RECT  4.735 0.495 4.825 1.185 ;
        RECT  4.625 0.495 4.735 0.600 ;
        RECT  4.645 1.060 4.735 1.185 ;
        RECT  3.775 1.195 4.355 1.325 ;
        RECT  3.775 0.475 4.345 0.585 ;
        RECT  3.670 0.475 3.775 1.325 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.370 1.255 3.460 1.525 ;
        RECT  3.330 1.075 3.440 1.165 ;
        RECT  1.530 1.255 3.370 1.345 ;
        RECT  2.995 0.475 3.340 0.585 ;
        RECT  3.160 0.255 3.330 0.365 ;
        RECT  2.995 1.055 3.220 1.165 ;
        RECT  1.670 0.275 3.160 0.365 ;
        RECT  2.905 0.475 2.995 1.165 ;
        RECT  2.595 0.475 2.905 0.585 ;
        RECT  2.555 1.055 2.905 1.165 ;
        RECT  1.750 0.475 2.305 0.580 ;
        RECT  1.750 1.055 2.265 1.165 ;
        RECT  1.640 0.475 1.750 1.165 ;
        RECT  1.460 0.255 1.670 0.365 ;
        RECT  1.530 0.475 1.545 0.565 ;
        RECT  1.440 0.475 1.530 1.345 ;
        RECT  0.195 0.275 1.460 0.365 ;
        RECT  1.375 0.475 1.440 0.565 ;
        RECT  1.435 1.075 1.440 1.345 ;
        RECT  1.300 1.075 1.435 1.165 ;
        RECT  1.050 0.475 1.285 0.565 ;
        RECT  1.050 1.075 1.190 1.165 ;
        RECT  0.195 1.435 1.120 1.525 ;
        RECT  0.960 0.475 1.050 1.165 ;
        RECT  0.740 0.475 0.960 0.565 ;
        RECT  0.545 1.075 0.960 1.165 ;
        RECT  0.650 0.475 0.740 0.645 ;
        RECT  0.140 0.275 0.195 0.560 ;
        RECT  0.140 1.220 0.195 1.525 ;
        RECT  0.050 0.275 0.140 1.525 ;
    END
END MUX4D4

MACRO MUX4ND0
    CLASS CORE ;
    FOREIGN MUX4ND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.890 0.710 3.950 1.135 ;
        RECT  3.850 0.710 3.890 1.345 ;
        RECT  3.840 0.710 3.850 0.820 ;
        RECT  3.790 1.025 3.850 1.345 ;
        RECT  3.730 0.440 3.840 0.820 ;
        RECT  3.700 1.235 3.790 1.345 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 0.710 3.155 1.090 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0836 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.710 1.750 1.090 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0326 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.090 ;
        RECT  1.095 0.710 1.250 0.925 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.950 1.090 ;
        RECT  2.775 0.710 2.850 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0331 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 1.965 1.090 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.165 4.200 0.165 ;
        RECT  1.655 -0.165 1.765 0.395 ;
        RECT  1.430 -0.165 1.655 0.165 ;
        RECT  1.320 -0.165 1.430 0.395 ;
        RECT  0.185 -0.165 1.320 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.635 4.200 1.965 ;
        RECT  1.670 1.445 1.880 1.965 ;
        RECT  1.330 1.635 1.670 1.965 ;
        RECT  1.120 1.445 1.330 1.965 ;
        RECT  0.185 1.635 1.120 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.060 0.485 4.150 1.525 ;
        RECT  3.940 0.485 4.060 0.595 ;
        RECT  3.990 1.245 4.060 1.525 ;
        RECT  2.170 1.435 3.990 1.525 ;
        RECT  3.510 0.275 3.610 1.345 ;
        RECT  3.470 0.275 3.510 0.650 ;
        RECT  3.440 1.235 3.510 1.345 ;
        RECT  2.455 0.275 3.470 0.365 ;
        RECT  3.355 0.880 3.420 1.090 ;
        RECT  3.350 0.490 3.355 1.090 ;
        RECT  3.260 0.490 3.350 1.345 ;
        RECT  3.155 0.490 3.260 0.600 ;
        RECT  3.155 1.235 3.260 1.345 ;
        RECT  2.655 0.475 2.780 0.585 ;
        RECT  2.655 1.200 2.755 1.310 ;
        RECT  2.545 0.475 2.655 1.310 ;
        RECT  2.345 0.275 2.455 1.320 ;
        RECT  1.945 0.315 2.245 0.425 ;
        RECT  2.060 1.265 2.170 1.525 ;
        RECT  2.055 0.515 2.165 1.175 ;
        RECT  0.725 1.265 2.060 1.355 ;
        RECT  1.855 0.315 1.945 0.600 ;
        RECT  1.535 0.505 1.855 0.600 ;
        RECT  1.440 0.505 1.535 1.155 ;
        RECT  1.195 0.505 1.440 0.615 ;
        RECT  1.095 0.315 1.195 0.615 ;
        RECT  0.730 0.315 1.095 0.425 ;
        RECT  0.880 0.515 0.990 1.175 ;
        RECT  0.605 0.515 0.725 1.355 ;
        RECT  0.335 0.280 0.445 1.365 ;
    END
END MUX4ND0

MACRO MUX4ND1
    CLASS CORE ;
    FOREIGN MUX4ND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.275 5.150 1.525 ;
        RECT  5.025 0.275 5.050 0.675 ;
        RECT  5.025 1.045 5.050 1.525 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0696 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.445 0.705 3.555 1.120 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.1070 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.710 1.755 1.120 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.120 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0327 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.120 ;
        RECT  1.095 0.710 1.245 0.925 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0555 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.705 2.955 1.120 ;
        RECT  2.775 0.705 2.845 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0326 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.710 1.965 1.120 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.165 5.200 0.165 ;
        RECT  1.655 -0.165 1.765 0.395 ;
        RECT  1.430 -0.165 1.655 0.165 ;
        RECT  1.320 -0.165 1.430 0.395 ;
        RECT  0.195 -0.165 1.320 0.165 ;
        RECT  0.065 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.635 5.200 1.965 ;
        RECT  1.690 1.445 1.860 1.965 ;
        RECT  1.305 1.635 1.690 1.965 ;
        RECT  1.135 1.445 1.305 1.965 ;
        RECT  0.195 1.635 1.135 1.965 ;
        RECT  0.065 1.240 0.195 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.915 0.750 4.960 0.920 ;
        RECT  4.825 0.275 4.915 0.920 ;
        RECT  4.255 0.275 4.825 0.365 ;
        RECT  4.710 1.025 4.800 1.525 ;
        RECT  4.700 0.740 4.710 1.525 ;
        RECT  4.620 0.740 4.700 1.125 ;
        RECT  2.170 1.435 4.700 1.525 ;
        RECT  4.505 1.215 4.610 1.325 ;
        RECT  4.505 0.475 4.590 0.605 ;
        RECT  4.395 0.475 4.505 1.325 ;
        RECT  4.255 1.235 4.285 1.345 ;
        RECT  4.145 0.275 4.255 1.345 ;
        RECT  4.115 1.235 4.145 1.345 ;
        RECT  4.000 1.235 4.025 1.345 ;
        RECT  3.900 0.275 4.000 1.345 ;
        RECT  3.880 0.275 3.900 0.675 ;
        RECT  3.855 1.235 3.900 1.345 ;
        RECT  3.315 0.275 3.880 0.365 ;
        RECT  3.770 0.890 3.805 1.080 ;
        RECT  3.765 0.475 3.770 1.080 ;
        RECT  3.675 0.475 3.765 1.345 ;
        RECT  3.580 0.475 3.675 0.585 ;
        RECT  3.585 1.235 3.675 1.345 ;
        RECT  3.225 0.275 3.315 1.320 ;
        RECT  3.100 0.275 3.225 0.415 ;
        RECT  3.100 1.140 3.225 1.320 ;
        RECT  3.045 0.525 3.135 0.930 ;
        RECT  2.950 0.525 3.045 0.615 ;
        RECT  2.860 0.275 2.950 0.615 ;
        RECT  2.455 0.275 2.860 0.365 ;
        RECT  2.655 0.475 2.770 0.585 ;
        RECT  2.655 1.140 2.745 1.320 ;
        RECT  2.545 0.475 2.655 1.320 ;
        RECT  2.345 0.275 2.455 1.320 ;
        RECT  1.945 0.315 2.255 0.425 ;
        RECT  2.060 1.265 2.170 1.525 ;
        RECT  2.055 0.515 2.165 1.175 ;
        RECT  0.725 1.265 2.060 1.355 ;
        RECT  1.855 0.315 1.945 0.600 ;
        RECT  1.535 0.505 1.855 0.600 ;
        RECT  1.445 0.505 1.535 1.155 ;
        RECT  1.195 0.505 1.445 0.615 ;
        RECT  1.095 0.315 1.195 0.615 ;
        RECT  0.730 0.315 1.095 0.425 ;
        RECT  0.875 0.515 0.985 1.175 ;
        RECT  0.605 0.515 0.725 1.355 ;
        RECT  0.335 0.275 0.445 1.355 ;
    END
END MUX4ND1

MACRO MUX4ND2
    CLASS CORE ;
    FOREIGN MUX4ND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.060 0.275 5.150 1.185 ;
        RECT  5.050 0.275 5.060 1.490 ;
        RECT  4.915 0.275 5.050 0.430 ;
        RECT  4.960 1.045 5.050 1.490 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0684 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.445 0.705 3.555 1.120 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.1069 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.710 1.755 1.120 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.120 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0327 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.355 1.120 ;
        RECT  1.095 0.710 1.245 0.925 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.705 2.955 1.120 ;
        RECT  2.775 0.705 2.845 0.920 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0326 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.710 1.965 1.120 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.165 5.400 0.165 ;
        RECT  1.655 -0.165 1.765 0.395 ;
        RECT  1.430 -0.165 1.655 0.165 ;
        RECT  1.320 -0.165 1.430 0.395 ;
        RECT  0.195 -0.165 1.320 0.165 ;
        RECT  0.065 -0.165 0.195 0.465 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.335 1.635 5.400 1.965 ;
        RECT  5.205 1.305 5.335 1.965 ;
        RECT  1.860 1.635 5.205 1.965 ;
        RECT  1.690 1.445 1.860 1.965 ;
        RECT  1.305 1.635 1.690 1.965 ;
        RECT  1.135 1.445 1.305 1.965 ;
        RECT  0.195 1.635 1.135 1.965 ;
        RECT  0.065 1.230 0.195 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.860 0.540 4.960 0.920 ;
        RECT  4.805 0.540 4.860 0.630 ;
        RECT  4.710 1.025 4.810 1.525 ;
        RECT  4.705 0.275 4.805 0.630 ;
        RECT  4.705 1.025 4.710 1.125 ;
        RECT  2.170 1.435 4.710 1.525 ;
        RECT  4.255 0.275 4.705 0.365 ;
        RECT  4.605 0.740 4.705 1.125 ;
        RECT  4.515 0.475 4.595 0.605 ;
        RECT  4.515 1.235 4.595 1.345 ;
        RECT  4.405 0.475 4.515 1.345 ;
        RECT  4.255 1.235 4.285 1.345 ;
        RECT  4.145 0.275 4.255 1.345 ;
        RECT  4.115 1.235 4.145 1.345 ;
        RECT  4.000 1.235 4.025 1.345 ;
        RECT  3.895 0.275 4.000 1.345 ;
        RECT  3.315 0.275 3.895 0.365 ;
        RECT  3.855 1.235 3.895 1.345 ;
        RECT  3.765 0.890 3.805 1.080 ;
        RECT  3.675 0.475 3.765 1.345 ;
        RECT  3.585 0.475 3.675 0.585 ;
        RECT  3.585 1.235 3.675 1.345 ;
        RECT  3.225 0.275 3.315 1.320 ;
        RECT  3.100 0.275 3.225 0.415 ;
        RECT  3.100 1.140 3.225 1.320 ;
        RECT  3.045 0.525 3.135 0.930 ;
        RECT  2.990 0.525 3.045 0.615 ;
        RECT  2.900 0.275 2.990 0.615 ;
        RECT  2.455 0.275 2.900 0.365 ;
        RECT  2.655 0.475 2.790 0.585 ;
        RECT  2.655 1.140 2.745 1.320 ;
        RECT  2.545 0.475 2.655 1.320 ;
        RECT  2.355 0.275 2.455 1.320 ;
        RECT  2.345 0.790 2.355 1.320 ;
        RECT  1.945 0.315 2.265 0.425 ;
        RECT  2.060 1.265 2.170 1.525 ;
        RECT  2.055 0.515 2.165 1.175 ;
        RECT  0.725 1.265 2.060 1.355 ;
        RECT  1.855 0.315 1.945 0.600 ;
        RECT  1.535 0.505 1.855 0.600 ;
        RECT  1.445 0.505 1.535 1.155 ;
        RECT  1.195 0.505 1.445 0.615 ;
        RECT  0.875 0.515 0.985 1.175 ;
        RECT  0.605 0.515 0.725 1.355 ;
        RECT  0.335 0.275 0.445 1.355 ;
        RECT  1.095 0.315 1.195 0.615 ;
        RECT  0.730 0.315 1.095 0.425 ;
    END
END MUX4ND2

MACRO MUX4ND4
    CLASS CORE ;
    FOREIGN MUX4ND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 0.310 8.105 0.690 ;
        RECT  8.050 1.110 8.105 1.490 ;
        RECT  7.750 0.310 8.050 1.490 ;
        RECT  7.415 0.310 7.750 0.690 ;
        RECT  7.415 1.110 7.750 1.490 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0941 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.445 0.680 5.555 1.120 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.1087 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.505 2.555 0.920 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.555 0.890 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0655 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.710 1.755 0.890 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.1106 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.710 4.355 0.925 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0625 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.710 3.155 0.905 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.335 -0.165 8.400 0.165 ;
        RECT  8.215 -0.165 8.335 0.690 ;
        RECT  3.105 -0.165 8.215 0.165 ;
        RECT  3.015 -0.165 3.105 0.395 ;
        RECT  1.640 -0.165 3.015 0.165 ;
        RECT  1.550 -0.165 1.640 0.395 ;
        RECT  0.455 -0.165 1.550 0.165 ;
        RECT  0.325 -0.165 0.455 0.535 ;
        RECT  0.000 -0.165 0.325 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.335 1.635 8.400 1.965 ;
        RECT  8.215 1.110 8.335 1.965 ;
        RECT  4.260 1.635 8.215 1.965 ;
        RECT  4.090 1.515 4.260 1.965 ;
        RECT  3.040 1.635 4.090 1.965 ;
        RECT  2.870 1.445 3.040 1.965 ;
        RECT  2.490 1.635 2.870 1.965 ;
        RECT  2.305 1.445 2.490 1.965 ;
        RECT  1.615 1.635 2.305 1.965 ;
        RECT  1.445 1.445 1.615 1.965 ;
        RECT  0.455 1.635 1.445 1.965 ;
        RECT  0.325 1.220 0.455 1.965 ;
        RECT  0.000 1.635 0.325 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.415 0.310 7.650 0.690 ;
        RECT  7.415 1.110 7.650 1.490 ;
        RECT  7.225 0.275 7.325 0.945 ;
        RECT  6.315 0.275 7.225 0.365 ;
        RECT  6.985 0.455 7.085 1.490 ;
        RECT  6.585 0.455 6.985 0.565 ;
        RECT  6.725 0.740 6.825 1.525 ;
        RECT  5.755 1.435 6.725 1.525 ;
        RECT  6.475 0.455 6.585 1.315 ;
        RECT  6.315 1.235 6.345 1.345 ;
        RECT  6.205 0.275 6.315 1.345 ;
        RECT  6.175 1.235 6.205 1.345 ;
        RECT  5.955 0.275 6.065 1.345 ;
        RECT  5.315 0.275 5.955 0.365 ;
        RECT  5.890 1.235 5.955 1.345 ;
        RECT  5.795 0.765 5.865 0.955 ;
        RECT  5.775 0.475 5.795 0.955 ;
        RECT  5.685 0.475 5.775 1.225 ;
        RECT  5.655 1.335 5.755 1.525 ;
        RECT  5.655 0.765 5.685 1.225 ;
        RECT  3.960 1.335 5.655 1.425 ;
        RECT  5.195 0.275 5.315 1.235 ;
        RECT  4.780 1.125 5.195 1.235 ;
        RECT  4.975 0.275 5.085 0.955 ;
        RECT  3.755 0.275 4.975 0.365 ;
        RECT  4.780 0.475 4.850 0.600 ;
        RECT  4.670 0.475 4.780 1.235 ;
        RECT  3.955 0.475 4.580 0.600 ;
        RECT  3.955 1.125 4.555 1.235 ;
        RECT  3.870 1.335 3.960 1.525 ;
        RECT  3.845 0.475 3.955 1.235 ;
        RECT  3.265 1.435 3.870 1.525 ;
        RECT  3.665 0.275 3.755 1.325 ;
        RECT  3.455 1.215 3.665 1.325 ;
        RECT  3.285 0.315 3.575 0.425 ;
        RECT  3.375 0.515 3.485 1.105 ;
        RECT  3.335 1.015 3.375 1.105 ;
        RECT  3.165 1.015 3.335 1.175 ;
        RECT  3.195 0.315 3.285 0.595 ;
        RECT  3.175 1.265 3.265 1.525 ;
        RECT  2.925 0.505 3.195 0.595 ;
        RECT  0.975 1.265 3.175 1.355 ;
        RECT  2.745 1.065 3.165 1.175 ;
        RECT  2.835 0.315 2.925 0.595 ;
        RECT  2.260 0.315 2.835 0.405 ;
        RECT  2.645 0.515 2.745 1.175 ;
        RECT  2.565 1.065 2.645 1.175 ;
        RECT  2.170 0.315 2.260 1.175 ;
        RECT  1.820 0.315 2.170 0.405 ;
        RECT  2.025 1.065 2.170 1.175 ;
        RECT  1.935 0.515 2.000 0.800 ;
        RECT  1.910 0.515 1.935 1.155 ;
        RECT  1.845 0.710 1.910 1.155 ;
        RECT  1.220 1.025 1.845 1.155 ;
        RECT  1.730 0.315 1.820 0.595 ;
        RECT  1.460 0.505 1.730 0.595 ;
        RECT  1.370 0.325 1.460 0.595 ;
        RECT  1.000 0.325 1.370 0.415 ;
        RECT  1.220 0.535 1.280 0.670 ;
        RECT  1.110 0.535 1.220 1.155 ;
        RECT  0.975 0.535 1.020 0.670 ;
        RECT  0.845 0.535 0.975 1.515 ;
        RECT  0.715 0.285 0.735 1.090 ;
        RECT  0.645 0.285 0.715 1.515 ;
        RECT  0.560 0.285 0.645 0.495 ;
        RECT  0.585 1.000 0.645 1.515 ;
        RECT  0.195 1.000 0.585 1.090 ;
        RECT  0.155 0.285 0.195 0.600 ;
        RECT  0.155 1.000 0.195 1.505 ;
        RECT  0.065 0.285 0.155 1.505 ;
    END
END MUX4ND4

MACRO ND2D0
    CLASS CORE ;
    FOREIGN ND2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.295 0.750 1.120 ;
        RECT  0.555 0.295 0.650 0.400 ;
        RECT  0.455 1.030 0.650 1.120 ;
        RECT  0.345 1.030 0.455 1.520 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.680 0.190 0.930 ;
        RECT  0.050 0.680 0.150 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.550 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.165 0.800 0.165 ;
        RECT  0.085 -0.165 0.195 0.460 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.230 0.715 1.965 ;
        RECT  0.195 1.635 0.605 1.965 ;
        RECT  0.085 1.230 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END ND2D0

MACRO ND2D1
    CLASS CORE ;
    FOREIGN ND2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.295 0.750 1.120 ;
        RECT  0.555 0.295 0.650 0.400 ;
        RECT  0.455 1.030 0.650 1.120 ;
        RECT  0.345 1.030 0.455 1.520 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.680 0.190 0.930 ;
        RECT  0.050 0.680 0.150 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.550 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.165 0.800 0.165 ;
        RECT  0.085 -0.165 0.195 0.560 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.635 0.800 1.965 ;
        RECT  0.605 1.230 0.715 1.965 ;
        RECT  0.195 1.635 0.605 1.965 ;
        RECT  0.085 1.230 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END ND2D1

MACRO ND2D2
    CLASS CORE ;
    FOREIGN ND2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 1.065 1.255 ;
        RECT  0.550 0.460 0.805 0.570 ;
        RECT  0.450 0.460 0.550 1.255 ;
        RECT  0.355 1.145 0.450 1.255 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.785 1.350 1.490 ;
        RECT  1.060 0.785 1.250 0.890 ;
        RECT  0.150 1.400 1.250 1.490 ;
        RECT  0.150 0.780 0.340 0.890 ;
        RECT  0.050 0.710 0.150 1.490 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 -0.165 1.400 0.165 ;
        RECT  1.165 -0.165 1.275 0.695 ;
        RECT  0.235 -0.165 1.165 0.165 ;
        RECT  0.125 -0.165 0.235 0.585 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.400 1.965 ;
        END
    END VDD
END ND2D2

MACRO ND2D3
    CLASS CORE ;
    FOREIGN ND2D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.635 0.350 1.725 1.140 ;
        RECT  1.615 0.350 1.635 0.595 ;
        RECT  1.460 1.050 1.635 1.140 ;
        RECT  0.545 0.350 1.615 0.460 ;
        RECT  1.150 1.050 1.460 1.350 ;
        RECT  0.285 1.180 1.150 1.275 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1651 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.780 1.265 0.890 ;
        RECT  0.895 0.780 0.995 1.090 ;
        RECT  0.350 1.000 0.895 1.090 ;
        RECT  0.250 0.680 0.350 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.525 0.730 1.545 0.940 ;
        RECT  1.435 0.570 1.525 0.940 ;
        RECT  0.750 0.570 1.435 0.660 ;
        RECT  0.655 0.570 0.750 0.890 ;
        RECT  0.450 0.710 0.655 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 1.800 0.165 ;
        RECT  0.075 -0.165 0.185 0.500 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.250 1.725 1.965 ;
        RECT  0.655 1.635 1.615 1.965 ;
        RECT  0.655 1.385 0.755 1.495 ;
        RECT  0.545 1.385 0.655 1.965 ;
        RECT  0.185 1.635 0.545 1.965 ;
        RECT  0.075 1.355 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.635 0.350 1.725 1.140 ;
        RECT  1.615 0.350 1.635 0.595 ;
        RECT  1.550 1.050 1.635 1.140 ;
        RECT  0.545 0.350 1.615 0.460 ;
        RECT  0.285 1.180 1.050 1.275 ;
    END
END ND2D3

MACRO ND2D4
    CLASS CORE ;
    FOREIGN ND2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 1.050 2.250 1.350 ;
        RECT  1.890 1.050 1.950 1.270 ;
        RECT  1.800 0.530 1.890 1.270 ;
        RECT  1.585 0.530 1.800 0.640 ;
        RECT  0.560 1.180 1.800 1.270 ;
        RECT  0.560 0.530 0.750 0.640 ;
        RECT  0.450 0.530 0.560 1.270 ;
        RECT  0.445 1.060 0.450 1.270 ;
        RECT  0.335 1.060 0.445 1.490 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2186 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 0.780 2.230 0.895 ;
        RECT  1.980 0.305 2.070 0.895 ;
        RECT  1.475 0.305 1.980 0.395 ;
        RECT  1.385 0.305 1.475 0.600 ;
        RECT  1.150 0.510 1.385 0.600 ;
        RECT  1.050 0.510 1.150 0.890 ;
        RECT  0.955 0.510 1.050 0.600 ;
        RECT  0.865 0.305 0.955 0.600 ;
        RECT  0.360 0.305 0.865 0.395 ;
        RECT  0.270 0.305 0.360 0.890 ;
        RECT  0.110 0.780 0.270 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.780 1.710 0.890 ;
        RECT  1.450 0.780 1.550 1.090 ;
        RECT  0.950 1.000 1.450 1.090 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.650 0.775 0.850 0.895 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 -0.165 2.400 0.165 ;
        RECT  2.180 -0.165 2.290 0.665 ;
        RECT  1.275 -0.165 2.180 0.165 ;
        RECT  1.065 -0.165 1.275 0.415 ;
        RECT  0.180 -0.165 1.065 0.165 ;
        RECT  0.070 -0.165 0.180 0.665 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.340 1.635 2.400 1.965 ;
        RECT  2.130 1.495 2.340 1.965 ;
        RECT  1.175 1.635 2.130 1.965 ;
        RECT  1.175 1.380 1.795 1.490 ;
        RECT  1.030 1.380 1.175 1.965 ;
        RECT  0.545 1.380 1.030 1.490 ;
        RECT  0.185 1.635 1.030 1.965 ;
        RECT  0.075 1.055 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END ND2D4

MACRO ND2D8
    CLASS CORE ;
    FOREIGN ND2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.1280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.900 1.180 4.115 1.290 ;
        RECT  3.800 0.510 3.900 1.290 ;
        RECT  3.575 0.510 3.800 0.620 ;
        RECT  2.665 1.180 3.800 1.290 ;
        RECT  2.665 0.510 2.835 0.620 ;
        RECT  2.575 0.510 2.665 1.290 ;
        RECT  2.450 1.180 2.575 1.290 ;
        RECT  2.150 1.050 2.450 1.350 ;
        RECT  1.845 1.180 2.150 1.290 ;
        RECT  1.755 0.510 1.845 1.290 ;
        RECT  1.585 0.510 1.755 0.620 ;
        RECT  0.540 1.180 1.755 1.290 ;
        RECT  0.540 0.510 0.740 0.620 ;
        RECT  0.450 0.510 0.540 1.290 ;
        RECT  0.285 1.180 0.450 1.290 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4189 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.105 0.785 4.245 0.890 ;
        RECT  4.015 0.310 4.105 0.890 ;
        RECT  3.355 0.310 4.015 0.400 ;
        RECT  3.245 0.310 3.355 0.910 ;
        RECT  2.465 0.310 3.245 0.400 ;
        RECT  2.375 0.310 2.465 0.890 ;
        RECT  2.045 0.780 2.375 0.890 ;
        RECT  1.955 0.310 2.045 0.890 ;
        RECT  1.475 0.310 1.955 0.400 ;
        RECT  1.385 0.310 1.475 0.600 ;
        RECT  1.350 0.510 1.385 0.600 ;
        RECT  1.235 0.510 1.350 0.890 ;
        RECT  0.955 0.510 1.235 0.600 ;
        RECT  1.160 0.780 1.235 0.890 ;
        RECT  0.850 0.310 0.955 0.600 ;
        RECT  0.360 0.310 0.850 0.400 ;
        RECT  0.270 0.310 0.360 0.890 ;
        RECT  0.110 0.785 0.270 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4183 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.710 1.645 0.940 ;
        RECT  1.450 0.710 1.550 1.090 ;
        RECT  0.765 1.000 1.450 1.090 ;
        RECT  0.650 0.710 0.765 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.675 ;
        RECT  2.265 -0.165 4.215 0.165 ;
        RECT  2.155 -0.165 2.265 0.665 ;
        RECT  1.175 -0.165 2.155 0.165 ;
        RECT  1.175 0.305 1.275 0.415 ;
        RECT  1.065 -0.165 1.175 0.415 ;
        RECT  0.180 -0.165 1.065 0.165 ;
        RECT  0.070 -0.165 0.180 0.675 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.090 4.325 1.965 ;
        RECT  3.370 1.635 4.215 1.965 ;
        RECT  3.370 1.380 3.855 1.490 ;
        RECT  3.230 1.380 3.370 1.965 ;
        RECT  2.605 1.380 3.230 1.490 ;
        RECT  1.170 1.635 3.230 1.965 ;
        RECT  1.170 1.380 1.795 1.490 ;
        RECT  1.030 1.380 1.170 1.965 ;
        RECT  0.545 1.380 1.030 1.490 ;
        RECT  0.185 1.635 1.030 1.965 ;
        RECT  0.075 1.045 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.900 1.180 4.115 1.290 ;
        RECT  3.800 0.510 3.900 1.290 ;
        RECT  3.575 0.510 3.800 0.620 ;
        RECT  2.665 1.180 3.800 1.290 ;
        RECT  2.665 0.510 2.835 0.620 ;
        RECT  2.575 0.510 2.665 1.290 ;
        RECT  2.550 1.180 2.575 1.290 ;
        RECT  1.845 1.180 2.050 1.290 ;
        RECT  1.755 0.510 1.845 1.290 ;
        RECT  1.585 0.510 1.755 0.620 ;
        RECT  0.540 1.180 1.755 1.290 ;
        RECT  0.540 0.510 0.740 0.620 ;
        RECT  0.450 0.510 0.540 1.290 ;
        RECT  0.285 1.180 0.450 1.290 ;
        RECT  3.570 0.730 3.680 1.090 ;
        RECT  2.880 1.000 3.570 1.090 ;
        RECT  2.775 0.730 2.880 1.090 ;
    END
END ND2D8

MACRO ND3D0
    CLASS CORE ;
    FOREIGN ND3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.130 ;
        RECT  0.965 0.510 1.050 0.600 ;
        RECT  0.965 1.040 1.050 1.130 ;
        RECT  0.850 0.310 0.965 0.600 ;
        RECT  0.850 1.040 0.965 1.490 ;
        RECT  0.445 1.040 0.850 1.130 ;
        RECT  0.335 1.040 0.445 1.470 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.750 0.800 0.920 ;
        RECT  0.650 0.510 0.750 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 1.200 0.165 ;
        RECT  0.075 -0.165 0.185 0.525 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.635 1.200 1.965 ;
        RECT  0.595 1.305 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.260 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END ND3D0

MACRO ND3D1
    CLASS CORE ;
    FOREIGN ND3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2910 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.130 ;
        RECT  0.965 0.510 1.050 0.600 ;
        RECT  0.965 1.040 1.050 1.130 ;
        RECT  0.850 0.310 0.965 0.600 ;
        RECT  0.850 1.040 0.965 1.490 ;
        RECT  0.445 1.040 0.850 1.130 ;
        RECT  0.335 1.040 0.445 1.470 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.750 0.800 0.920 ;
        RECT  0.650 0.510 0.750 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 1.200 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.635 1.200 1.965 ;
        RECT  0.595 1.305 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END ND3D1

MACRO ND3D2
    CLASS CORE ;
    FOREIGN ND3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.480 1.750 1.300 ;
        RECT  1.470 0.480 1.650 0.570 ;
        RECT  0.285 1.200 1.650 1.300 ;
        RECT  1.380 0.310 1.470 0.570 ;
        RECT  0.785 0.310 1.380 0.420 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1099 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.550 1.090 ;
        RECT  0.350 1.000 1.450 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        RECT  0.165 0.710 0.250 0.940 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1098 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.780 1.350 0.890 ;
        RECT  1.050 0.510 1.150 0.890 ;
        RECT  0.550 0.510 1.050 0.600 ;
        RECT  0.450 0.510 0.550 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.690 -0.165 1.800 0.165 ;
        RECT  1.580 -0.165 1.690 0.355 ;
        RECT  0.185 -0.165 1.580 0.165 ;
        RECT  0.075 -0.165 0.185 0.570 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.255 1.635 1.800 1.965 ;
        RECT  1.045 1.390 1.255 1.965 ;
        RECT  0.185 1.635 1.045 1.965 ;
        RECT  0.075 1.230 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END ND3D2

MACRO ND3D3
    CLASS CORE ;
    FOREIGN ND3D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6390 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.460 0.375 2.550 1.220 ;
        RECT  2.415 0.375 2.460 0.585 ;
        RECT  2.450 1.050 2.460 1.220 ;
        RECT  2.150 1.050 2.450 1.475 ;
        RECT  0.360 1.380 2.150 1.475 ;
        RECT  0.385 0.305 0.995 0.415 ;
        RECT  0.295 0.305 0.385 0.645 ;
        RECT  0.270 1.155 0.360 1.475 ;
        RECT  0.150 0.555 0.295 0.645 ;
        RECT  0.150 1.155 0.270 1.245 ;
        RECT  0.050 0.555 0.150 1.245 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1651 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.770 1.760 1.290 ;
        RECT  0.560 1.200 1.650 1.290 ;
        RECT  0.470 0.955 0.560 1.290 ;
        RECT  0.360 0.955 0.470 1.045 ;
        RECT  0.260 0.755 0.360 1.045 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1645 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.565 2.100 0.925 ;
        RECT  1.550 0.565 1.990 0.655 ;
        RECT  1.450 0.565 1.550 0.890 ;
        RECT  1.350 0.710 1.450 0.890 ;
        RECT  1.250 0.710 1.350 1.090 ;
        RECT  0.750 1.000 1.250 1.090 ;
        RECT  0.650 0.755 0.750 1.090 ;
        RECT  0.470 0.755 0.650 0.865 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1649 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.305 0.710 2.370 0.925 ;
        RECT  2.215 0.385 2.305 0.925 ;
        RECT  1.350 0.385 2.215 0.475 ;
        RECT  1.250 0.385 1.350 0.600 ;
        RECT  1.150 0.510 1.250 0.600 ;
        RECT  1.050 0.510 1.150 0.690 ;
        RECT  0.940 0.510 1.050 0.875 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.165 2.600 0.165 ;
        RECT  1.580 -0.165 1.765 0.295 ;
        RECT  0.185 -0.165 1.580 0.165 ;
        RECT  0.075 -0.165 0.185 0.445 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 1.635 2.600 1.965 ;
        RECT  0.070 1.355 0.180 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.460 0.375 2.550 0.950 ;
        RECT  2.415 0.375 2.460 0.585 ;
        RECT  0.360 1.380 2.050 1.475 ;
        RECT  0.385 0.305 0.995 0.415 ;
        RECT  0.295 0.305 0.385 0.645 ;
        RECT  0.270 1.155 0.360 1.475 ;
        RECT  0.150 0.555 0.295 0.645 ;
        RECT  0.150 1.155 0.270 1.245 ;
        RECT  0.050 0.555 0.150 1.245 ;
    END
END ND3D3

MACRO ND3D4
    CLASS CORE ;
    FOREIGN ND3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.285 3.350 1.505 ;
        RECT  2.370 0.285 3.250 0.390 ;
        RECT  0.150 1.360 3.250 1.505 ;
        RECT  0.150 0.285 1.030 0.390 ;
        RECT  0.050 0.285 0.150 1.505 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.2197 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.020 0.480 3.150 0.920 ;
        RECT  1.750 0.480 3.020 0.570 ;
        RECT  1.650 0.480 1.750 0.890 ;
        RECT  0.350 0.480 1.650 0.570 ;
        RECT  0.240 0.480 0.350 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2182 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.775 0.750 2.905 1.270 ;
        RECT  2.195 1.180 2.775 1.270 ;
        RECT  2.025 0.840 2.195 1.270 ;
        RECT  1.375 1.180 2.025 1.270 ;
        RECT  1.205 0.840 1.375 1.270 ;
        RECT  0.550 1.180 1.205 1.270 ;
        RECT  0.550 0.710 0.615 0.920 ;
        RECT  0.450 0.710 0.550 1.270 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2182 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.660 2.550 1.090 ;
        RECT  1.935 0.660 2.440 0.750 ;
        RECT  1.845 0.660 1.935 1.090 ;
        RECT  1.555 1.000 1.845 1.090 ;
        RECT  1.465 0.660 1.555 1.090 ;
        RECT  0.955 0.660 1.465 0.750 ;
        RECT  0.850 0.660 0.955 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.165 3.400 0.165 ;
        RECT  1.600 -0.165 1.770 0.390 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 3.400 1.965 ;
        END
    END VDD
END ND3D4

MACRO ND3D8
    CLASS CORE ;
    FOREIGN ND3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.5600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 1.120 6.475 1.290 ;
        RECT  6.050 0.510 6.465 0.680 ;
        RECT  5.750 0.510 6.050 1.290 ;
        RECT  4.715 0.510 5.750 0.620 ;
        RECT  0.285 1.120 5.750 1.290 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.4391 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 1.605 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4391 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 3.605 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4391 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 5.610 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.165 6.800 0.165 ;
        RECT  1.770 0.310 2.055 0.420 ;
        RECT  1.630 -0.165 1.770 0.420 ;
        RECT  0.770 -0.165 1.630 0.165 ;
        RECT  1.325 0.310 1.630 0.420 ;
        RECT  0.770 0.310 1.015 0.420 ;
        RECT  0.630 -0.165 0.770 0.420 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.295 0.310 0.630 0.420 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.685 1.635 6.800 1.965 ;
        RECT  6.575 1.040 6.685 1.965 ;
        RECT  5.770 1.635 6.575 1.965 ;
        RECT  5.770 1.380 6.215 1.490 ;
        RECT  5.630 1.380 5.770 1.965 ;
        RECT  4.965 1.380 5.630 1.490 ;
        RECT  4.170 1.635 5.630 1.965 ;
        RECT  4.170 1.380 4.655 1.490 ;
        RECT  4.030 1.380 4.170 1.965 ;
        RECT  3.665 1.380 4.030 1.490 ;
        RECT  3.170 1.635 4.030 1.965 ;
        RECT  3.170 1.380 3.355 1.490 ;
        RECT  3.030 1.380 3.170 1.965 ;
        RECT  2.625 1.380 3.030 1.490 ;
        RECT  1.970 1.635 3.030 1.965 ;
        RECT  1.970 1.380 2.315 1.490 ;
        RECT  1.830 1.380 1.970 1.965 ;
        RECT  1.585 1.380 1.830 1.490 ;
        RECT  0.970 1.635 1.830 1.965 ;
        RECT  0.970 1.380 1.275 1.490 ;
        RECT  0.830 1.380 0.970 1.965 ;
        RECT  0.545 1.380 0.830 1.490 ;
        RECT  0.185 1.635 0.830 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.150 1.120 6.475 1.290 ;
        RECT  6.150 0.510 6.465 0.680 ;
        RECT  4.715 0.510 5.650 0.620 ;
        RECT  0.285 1.120 5.650 1.290 ;
        RECT  6.575 0.310 6.685 0.585 ;
        RECT  4.605 0.310 6.575 0.420 ;
        RECT  4.495 0.310 4.605 0.680 ;
        RECT  2.365 0.310 4.495 0.420 ;
        RECT  0.185 0.510 4.385 0.620 ;
        RECT  0.075 0.375 0.185 0.620 ;
    END
END ND3D8

MACRO ND4D0
    CLASS CORE ;
    FOREIGN ND4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1430 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.300 1.350 1.150 ;
        RECT  1.065 0.300 1.250 0.400 ;
        RECT  0.965 1.060 1.250 1.150 ;
        RECT  0.850 1.060 0.965 1.490 ;
        RECT  0.450 1.060 0.850 1.150 ;
        RECT  0.335 1.060 0.450 1.490 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.240 0.890 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.750 0.790 0.920 ;
        RECT  0.650 0.510 0.750 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.510 1.150 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 1.400 0.165 ;
        RECT  0.075 -0.165 0.185 0.475 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 1.635 1.400 1.965 ;
        RECT  1.115 1.260 1.225 1.965 ;
        RECT  0.705 1.635 1.115 1.965 ;
        RECT  0.595 1.260 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.260 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END ND4D0

MACRO ND4D1
    CLASS CORE ;
    FOREIGN ND4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.300 1.350 1.150 ;
        RECT  1.065 0.300 1.250 0.400 ;
        RECT  0.965 1.060 1.250 1.150 ;
        RECT  0.850 1.060 0.965 1.490 ;
        RECT  0.450 1.060 0.850 1.150 ;
        RECT  0.335 1.060 0.450 1.490 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.240 0.890 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.510 0.550 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.750 0.790 0.920 ;
        RECT  0.650 0.510 0.750 0.920 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.510 1.150 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 1.400 0.165 ;
        RECT  0.075 -0.165 0.185 0.570 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 1.635 1.400 1.965 ;
        RECT  1.115 1.260 1.225 1.965 ;
        RECT  0.705 1.635 1.115 1.965 ;
        RECT  0.595 1.260 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.260 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END ND4D1

MACRO ND4D2
    CLASS CORE ;
    FOREIGN ND4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4940 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 1.035 2.265 1.490 ;
        RECT  1.750 1.035 2.155 1.125 ;
        RECT  1.635 1.035 1.750 1.490 ;
        RECT  0.965 1.035 1.635 1.125 ;
        RECT  0.850 1.035 0.965 1.490 ;
        RECT  0.550 1.035 0.850 1.125 ;
        RECT  0.450 0.500 0.550 1.125 ;
        RECT  0.295 0.500 0.450 0.600 ;
        RECT  0.445 1.035 0.450 1.125 ;
        RECT  0.335 1.035 0.445 1.490 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.350 0.890 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 1.150 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.340 0.890 ;
        RECT  0.050 0.680 0.150 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.215 -0.165 2.600 0.165 ;
        RECT  2.215 0.310 2.305 0.420 ;
        RECT  2.125 -0.165 2.215 0.420 ;
        RECT  0.000 -0.165 2.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.525 1.635 2.600 1.965 ;
        RECT  2.415 1.040 2.525 1.965 ;
        RECT  2.010 1.635 2.415 1.965 ;
        RECT  1.890 1.235 2.010 1.965 ;
        RECT  1.485 1.635 1.890 1.965 ;
        RECT  1.370 1.235 1.485 1.965 ;
        RECT  1.225 1.635 1.370 1.965 ;
        RECT  1.115 1.235 1.225 1.965 ;
        RECT  0.705 1.635 1.115 1.965 ;
        RECT  0.595 1.235 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.275 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.415 0.410 2.525 0.620 ;
        RECT  2.035 0.530 2.415 0.620 ;
        RECT  1.945 0.305 2.035 0.620 ;
        RECT  1.345 0.305 1.945 0.410 ;
        RECT  0.805 0.520 1.795 0.620 ;
        RECT  0.185 0.305 1.255 0.410 ;
        RECT  0.075 0.305 0.185 0.515 ;
    END
END ND4D2

MACRO ND4D3
    CLASS CORE ;
    FOREIGN ND4D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8370 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.195 1.035 3.350 1.505 ;
        RECT  2.785 1.035 3.195 1.165 ;
        RECT  2.650 1.035 2.785 1.505 ;
        RECT  2.265 1.035 2.650 1.165 ;
        RECT  2.155 1.035 2.265 1.505 ;
        RECT  1.750 1.035 2.155 1.165 ;
        RECT  1.635 1.035 1.750 1.505 ;
        RECT  1.225 1.035 1.635 1.165 ;
        RECT  1.115 1.035 1.225 1.505 ;
        RECT  0.850 1.035 1.115 1.165 ;
        RECT  0.750 0.500 0.850 1.165 ;
        RECT  0.595 0.500 0.750 1.505 ;
        RECT  0.550 0.500 0.595 1.165 ;
        RECT  0.185 0.500 0.550 0.600 ;
        RECT  0.185 1.035 0.550 1.165 ;
        RECT  0.075 0.310 0.185 0.600 ;
        RECT  0.050 1.035 0.185 1.505 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 3.150 0.890 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.350 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.550 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.430 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 -0.165 3.400 0.165 ;
        RECT  3.195 -0.165 3.305 0.585 ;
        RECT  2.970 -0.165 3.195 0.165 ;
        RECT  2.830 -0.165 2.970 0.420 ;
        RECT  0.000 -0.165 2.830 0.165 ;
        RECT  2.635 0.300 2.830 0.420 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.045 1.635 3.400 1.965 ;
        RECT  2.935 1.285 3.045 1.965 ;
        RECT  2.525 1.635 2.935 1.965 ;
        RECT  2.415 1.285 2.525 1.965 ;
        RECT  2.005 1.635 2.415 1.965 ;
        RECT  1.895 1.285 2.005 1.965 ;
        RECT  1.485 1.635 1.895 1.965 ;
        RECT  1.375 1.285 1.485 1.965 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.860 1.285 0.965 1.965 ;
        RECT  0.445 1.635 0.860 1.965 ;
        RECT  0.335 1.285 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.195 1.035 3.350 1.505 ;
        RECT  2.785 1.035 3.195 1.165 ;
        RECT  2.650 1.035 2.785 1.505 ;
        RECT  2.265 1.035 2.650 1.165 ;
        RECT  2.155 1.035 2.265 1.505 ;
        RECT  1.750 1.035 2.155 1.165 ;
        RECT  1.635 1.035 1.750 1.505 ;
        RECT  1.225 1.035 1.635 1.165 ;
        RECT  1.115 1.035 1.225 1.505 ;
        RECT  0.950 1.035 1.115 1.165 ;
        RECT  0.185 0.500 0.450 0.600 ;
        RECT  0.185 1.035 0.450 1.165 ;
        RECT  0.075 0.310 0.185 0.600 ;
        RECT  0.050 1.035 0.185 1.505 ;
        RECT  2.525 0.510 3.095 0.620 ;
        RECT  2.415 0.305 2.525 0.620 ;
        RECT  1.845 0.305 2.415 0.410 ;
        RECT  1.065 0.520 2.305 0.620 ;
        RECT  0.295 0.305 1.535 0.410 ;
    END
END ND4D3

MACRO ND4D4
    CLASS CORE ;
    FOREIGN ND4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.000 4.435 1.505 ;
        RECT  3.950 1.000 4.325 1.165 ;
        RECT  3.805 1.000 3.950 1.505 ;
        RECT  3.395 1.000 3.805 1.165 ;
        RECT  3.250 1.000 3.395 1.505 ;
        RECT  2.875 1.000 3.250 1.165 ;
        RECT  2.765 1.000 2.875 1.505 ;
        RECT  2.035 1.000 2.765 1.165 ;
        RECT  1.925 1.000 2.035 1.505 ;
        RECT  1.550 1.000 1.925 1.165 ;
        RECT  1.405 1.000 1.550 1.505 ;
        RECT  1.250 1.000 1.405 1.165 ;
        RECT  0.995 0.520 1.250 1.165 ;
        RECT  0.950 0.520 0.995 1.505 ;
        RECT  0.325 0.520 0.950 0.620 ;
        RECT  0.850 1.000 0.950 1.505 ;
        RECT  0.475 1.000 0.850 1.165 ;
        RECT  0.365 1.000 0.475 1.505 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.540 0.890 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.660 0.710 3.370 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 2.140 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.710 0.750 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 -0.165 4.800 0.165 ;
        RECT  4.170 0.310 4.485 0.420 ;
        RECT  4.030 -0.165 4.170 0.420 ;
        RECT  0.000 -0.165 4.030 0.165 ;
        RECT  3.755 0.310 4.030 0.420 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.695 1.635 4.800 1.965 ;
        RECT  4.585 1.045 4.695 1.965 ;
        RECT  4.175 1.635 4.585 1.965 ;
        RECT  4.065 1.285 4.175 1.965 ;
        RECT  3.655 1.635 4.065 1.965 ;
        RECT  3.545 1.285 3.655 1.965 ;
        RECT  3.135 1.635 3.545 1.965 ;
        RECT  3.025 1.285 3.135 1.965 ;
        RECT  2.615 1.635 3.025 1.965 ;
        RECT  2.505 1.285 2.615 1.965 ;
        RECT  2.295 1.635 2.505 1.965 ;
        RECT  2.185 1.285 2.295 1.965 ;
        RECT  1.775 1.635 2.185 1.965 ;
        RECT  1.665 1.285 1.775 1.965 ;
        RECT  1.255 1.635 1.665 1.965 ;
        RECT  1.145 1.285 1.255 1.965 ;
        RECT  0.735 1.635 1.145 1.965 ;
        RECT  0.625 1.285 0.735 1.965 ;
        RECT  0.215 1.635 0.625 1.965 ;
        RECT  0.105 1.045 0.215 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.325 1.000 4.435 1.505 ;
        RECT  3.950 1.000 4.325 1.165 ;
        RECT  3.805 1.000 3.950 1.505 ;
        RECT  3.395 1.000 3.805 1.165 ;
        RECT  3.250 1.000 3.395 1.505 ;
        RECT  2.875 1.000 3.250 1.165 ;
        RECT  2.765 1.000 2.875 1.505 ;
        RECT  2.035 1.000 2.765 1.165 ;
        RECT  1.925 1.000 2.035 1.505 ;
        RECT  1.550 1.000 1.925 1.165 ;
        RECT  1.405 1.000 1.550 1.505 ;
        RECT  1.350 1.000 1.405 1.165 ;
        RECT  0.325 0.520 0.850 0.620 ;
        RECT  0.475 1.000 0.850 1.165 ;
        RECT  0.365 1.000 0.475 1.505 ;
        RECT  4.585 0.375 4.695 0.620 ;
        RECT  3.655 0.530 4.585 0.620 ;
        RECT  3.545 0.305 3.655 0.620 ;
        RECT  2.455 0.305 3.545 0.410 ;
        RECT  1.365 0.520 3.435 0.620 ;
        RECT  0.215 0.305 2.345 0.410 ;
        RECT  0.105 0.305 0.215 0.585 ;
    END
END ND4D4

MACRO ND4D8
    CLASS CORE ;
    FOREIGN ND4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 3.105 0.680 ;
        RECT  2.250 1.015 3.105 1.115 ;
        RECT  1.950 0.510 2.250 1.115 ;
        RECT  1.335 0.510 1.950 0.680 ;
        RECT  1.355 1.015 1.950 1.115 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.165 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.780 0.710 0.850 0.930 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.670 0.550 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.835 -0.165 4.200 0.165 ;
        RECT  3.725 -0.165 3.835 0.495 ;
        RECT  3.315 -0.165 3.725 0.165 ;
        RECT  3.205 -0.165 3.315 0.495 ;
        RECT  2.570 -0.165 3.205 0.165 ;
        RECT  2.570 0.305 2.845 0.415 ;
        RECT  2.430 -0.165 2.570 0.415 ;
        RECT  1.570 -0.165 2.430 0.165 ;
        RECT  2.115 0.305 2.430 0.415 ;
        RECT  1.570 0.305 1.805 0.415 ;
        RECT  1.430 -0.165 1.570 0.415 ;
        RECT  0.000 -0.165 1.430 0.165 ;
        RECT  1.235 0.305 1.430 0.415 ;
        RECT  1.125 0.305 1.235 0.585 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.635 4.200 1.965 ;
        RECT  3.370 1.385 3.885 1.495 ;
        RECT  3.230 1.385 3.370 1.965 ;
        RECT  2.635 1.385 3.230 1.495 ;
        RECT  1.970 1.635 3.230 1.965 ;
        RECT  1.970 1.385 2.325 1.495 ;
        RECT  1.830 1.385 1.970 1.965 ;
        RECT  1.595 1.385 1.830 1.495 ;
        RECT  0.770 1.635 1.830 1.965 ;
        RECT  0.770 1.385 1.285 1.495 ;
        RECT  0.630 1.385 0.770 1.965 ;
        RECT  0.055 1.385 0.630 1.495 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.355 0.510 3.105 0.680 ;
        RECT  2.355 1.015 3.105 1.115 ;
        RECT  1.335 0.510 1.855 0.680 ;
        RECT  1.355 1.015 1.855 1.115 ;
        RECT  3.985 0.375 4.095 1.470 ;
        RECT  3.575 0.605 3.985 0.695 ;
        RECT  3.415 1.160 3.985 1.270 ;
        RECT  3.530 0.785 3.870 0.890 ;
        RECT  3.465 0.375 3.575 0.695 ;
        RECT  3.440 0.785 3.530 1.070 ;
        RECT  3.305 0.605 3.465 0.695 ;
        RECT  3.305 0.980 3.440 1.070 ;
        RECT  3.215 0.605 3.305 0.890 ;
        RECT  3.215 0.980 3.305 1.295 ;
        RECT  2.570 0.775 3.215 0.890 ;
        RECT  0.360 1.205 3.215 1.295 ;
        RECT  0.270 0.425 0.360 1.295 ;
        RECT  0.055 0.425 0.270 0.535 ;
    END
END ND4D8

MACRO NR2D0
    CLASS CORE ;
    FOREIGN NR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.510 0.750 1.340 ;
        RECT  0.455 0.510 0.650 0.600 ;
        RECT  0.555 1.230 0.650 1.340 ;
        RECT  0.345 0.280 0.455 0.600 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.240 0.890 ;
        RECT  0.050 0.680 0.150 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.655 -0.165 0.800 0.165 ;
        RECT  0.655 0.300 0.745 0.400 ;
        RECT  0.565 -0.165 0.655 0.400 ;
        RECT  0.195 -0.165 0.565 0.165 ;
        RECT  0.085 -0.165 0.195 0.475 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 1.635 0.800 1.965 ;
        RECT  0.085 1.240 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END NR2D0

MACRO NR2D1
    CLASS CORE ;
    FOREIGN NR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1660 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.510 0.750 1.340 ;
        RECT  0.455 0.510 0.650 0.600 ;
        RECT  0.555 1.230 0.650 1.340 ;
        RECT  0.345 0.280 0.455 0.600 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.240 0.890 ;
        RECT  0.050 0.680 0.150 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.655 -0.165 0.800 0.165 ;
        RECT  0.655 0.300 0.745 0.400 ;
        RECT  0.565 -0.165 0.655 0.400 ;
        RECT  0.195 -0.165 0.565 0.165 ;
        RECT  0.085 -0.165 0.195 0.570 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 1.635 0.800 1.965 ;
        RECT  0.085 1.240 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END NR2D1

MACRO NR2D2
    CLASS CORE ;
    FOREIGN NR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.905 0.310 1.015 0.600 ;
        RECT  0.555 0.510 0.905 0.600 ;
        RECT  0.555 1.205 0.805 1.315 ;
        RECT  0.495 0.510 0.555 1.315 ;
        RECT  0.445 0.310 0.495 1.315 ;
        RECT  0.385 0.310 0.445 0.600 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1108 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.710 1.155 1.205 ;
        RECT  1.045 0.710 1.135 1.515 ;
        RECT  0.355 1.425 1.045 1.515 ;
        RECT  0.265 0.710 0.355 1.515 ;
        RECT  0.245 0.710 0.265 1.205 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1104 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.710 0.755 1.095 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 -0.165 1.400 0.165 ;
        RECT  1.165 -0.165 1.275 0.540 ;
        RECT  0.805 -0.165 1.165 0.165 ;
        RECT  0.595 -0.165 0.805 0.400 ;
        RECT  0.235 -0.165 0.595 0.165 ;
        RECT  0.125 -0.165 0.235 0.540 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.335 1.635 1.400 1.965 ;
        RECT  1.225 1.315 1.335 1.965 ;
        RECT  0.175 1.635 1.225 1.965 ;
        RECT  0.075 1.315 0.175 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END NR2D2

MACRO NR2D3
    CLASS CORE ;
    FOREIGN NR2D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4210 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.375 1.750 1.350 ;
        RECT  0.285 0.375 1.650 0.485 ;
        RECT  1.350 1.050 1.650 1.350 ;
        RECT  0.545 1.240 1.350 1.350 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1651 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.795 1.270 0.900 ;
        RECT  1.050 0.795 1.150 1.120 ;
        RECT  0.350 1.030 1.050 1.120 ;
        RECT  0.250 0.680 0.350 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1651 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.595 1.550 0.940 ;
        RECT  0.950 0.595 1.450 0.685 ;
        RECT  0.850 0.595 0.950 0.890 ;
        RECT  0.650 0.710 0.850 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 1.800 0.165 ;
        RECT  0.075 -0.165 0.185 0.585 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.635 1.800 1.965 ;
        RECT  0.075 1.230 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.650 0.375 1.750 0.950 ;
        RECT  0.285 0.375 1.650 0.485 ;
        RECT  0.545 1.240 1.250 1.350 ;
    END
END NR2D3

MACRO NR2D4
    CLASS CORE ;
    FOREIGN NR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.895 0.325 2.085 0.475 ;
        RECT  1.805 0.325 1.895 1.295 ;
        RECT  1.550 0.325 1.805 0.745 ;
        RECT  1.615 1.125 1.805 1.295 ;
        RECT  0.550 0.325 1.550 0.485 ;
        RECT  0.550 1.200 0.805 1.310 ;
        RECT  0.450 0.325 0.550 1.310 ;
        RECT  0.335 0.325 0.450 0.485 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2197 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.765 2.120 1.515 ;
        RECT  1.155 1.420 2.010 1.515 ;
        RECT  1.045 0.775 1.155 1.515 ;
        RECT  0.360 1.420 1.045 1.515 ;
        RECT  0.270 0.770 0.360 1.515 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.835 1.695 0.935 ;
        RECT  1.285 0.595 1.375 0.935 ;
        RECT  0.755 0.595 1.285 0.685 ;
        RECT  0.645 0.595 0.755 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.305 -0.165 2.400 0.165 ;
        RECT  2.195 -0.165 2.305 0.675 ;
        RECT  0.235 -0.165 2.195 0.165 ;
        RECT  0.125 -0.165 0.235 0.675 ;
        RECT  0.000 -0.165 0.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.635 2.400 1.965 ;
        RECT  2.210 1.040 2.320 1.965 ;
        RECT  0.180 1.635 2.210 1.965 ;
        RECT  0.080 1.040 0.180 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.920 0.325 2.085 0.475 ;
        RECT  1.805 0.820 1.895 1.295 ;
        RECT  1.615 1.125 1.805 1.295 ;
        RECT  0.550 0.325 1.480 0.485 ;
        RECT  0.550 1.200 0.805 1.310 ;
        RECT  0.450 0.325 0.550 1.310 ;
        RECT  0.335 0.325 0.450 0.485 ;
    END
END NR2D4

MACRO NR2D8
    CLASS CORE ;
    FOREIGN NR2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.0400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.505 4.115 0.675 ;
        RECT  3.450 1.070 4.115 1.240 ;
        RECT  3.150 0.505 3.450 1.240 ;
        RECT  0.285 0.505 3.150 0.605 ;
        RECT  2.345 1.070 3.150 1.240 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4381 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 1.605 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 3.000 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.695 ;
        RECT  3.570 -0.165 4.215 0.165 ;
        RECT  3.570 0.305 3.855 0.415 ;
        RECT  3.430 -0.165 3.570 0.415 ;
        RECT  2.570 -0.165 3.430 0.165 ;
        RECT  3.125 0.305 3.430 0.415 ;
        RECT  2.570 0.305 2.815 0.415 ;
        RECT  2.430 -0.165 2.570 0.415 ;
        RECT  0.970 -0.165 2.430 0.165 ;
        RECT  2.085 0.305 2.430 0.415 ;
        RECT  0.970 0.305 1.275 0.415 ;
        RECT  0.830 -0.165 0.970 0.415 ;
        RECT  0.185 -0.165 0.830 0.165 ;
        RECT  0.545 0.305 0.830 0.415 ;
        RECT  0.075 -0.165 0.185 0.695 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 1.635 4.400 1.965 ;
        RECT  1.375 1.280 1.485 1.965 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.855 1.280 0.965 1.965 ;
        RECT  0.445 1.635 0.855 1.965 ;
        RECT  0.335 1.280 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.550 0.505 4.115 0.675 ;
        RECT  3.550 1.070 4.115 1.240 ;
        RECT  0.285 0.505 3.050 0.605 ;
        RECT  2.345 1.070 3.050 1.240 ;
        RECT  4.215 1.030 4.325 1.490 ;
        RECT  2.245 1.375 4.215 1.490 ;
        RECT  2.135 1.060 2.245 1.490 ;
        RECT  0.185 1.060 2.135 1.170 ;
        RECT  0.075 1.060 0.185 1.515 ;
    END
END NR2D8

MACRO NR2XD0
    CLASS CORE ;
    FOREIGN NR2XD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.510 0.750 1.340 ;
        RECT  0.455 0.510 0.650 0.600 ;
        RECT  0.555 1.230 0.650 1.340 ;
        RECT  0.345 0.280 0.455 0.600 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.780 0.240 0.890 ;
        RECT  0.050 0.680 0.150 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.655 -0.165 0.800 0.165 ;
        RECT  0.655 0.300 0.745 0.400 ;
        RECT  0.565 -0.165 0.655 0.400 ;
        RECT  0.195 -0.165 0.565 0.165 ;
        RECT  0.085 -0.165 0.195 0.475 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 1.635 0.800 1.965 ;
        RECT  0.085 1.240 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
END NR2XD0

MACRO NR2XD1
    CLASS CORE ;
    FOREIGN NR2XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 1.010 1.065 1.120 ;
        RECT  0.645 0.270 0.755 1.120 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 1.150 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.165 1.400 0.165 ;
        RECT  0.905 -0.165 1.015 0.580 ;
        RECT  0.495 -0.165 0.905 0.165 ;
        RECT  0.385 -0.165 0.495 0.580 ;
        RECT  0.000 -0.165 0.385 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.445 1.635 1.400 1.965 ;
        RECT  0.445 1.395 0.545 1.505 ;
        RECT  0.335 1.395 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.165 1.040 1.275 1.470 ;
        RECT  0.235 1.210 1.165 1.305 ;
        RECT  0.125 1.040 0.235 1.470 ;
    END
END NR2XD1

MACRO NR2XD2
    CLASS CORE ;
    FOREIGN NR2XD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.010 2.085 1.120 ;
        RECT  1.405 0.270 1.550 0.690 ;
        RECT  1.350 0.575 1.405 0.690 ;
        RECT  1.250 0.575 1.350 1.120 ;
        RECT  0.995 0.575 1.250 0.690 ;
        RECT  0.850 0.270 0.995 0.690 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1716 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.780 1.100 0.890 ;
        RECT  0.250 0.710 0.750 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1716 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 2.150 0.890 ;
        RECT  1.490 0.780 1.650 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.775 -0.165 2.400 0.165 ;
        RECT  1.665 -0.165 1.775 0.580 ;
        RECT  1.255 -0.165 1.665 0.165 ;
        RECT  1.145 -0.165 1.255 0.485 ;
        RECT  0.735 -0.165 1.145 0.165 ;
        RECT  0.625 -0.165 0.735 0.580 ;
        RECT  0.000 -0.165 0.625 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 1.635 2.400 1.965 ;
        RECT  0.945 1.395 1.045 1.505 ;
        RECT  0.835 1.395 0.945 1.965 ;
        RECT  0.475 1.635 0.835 1.965 ;
        RECT  0.365 1.240 0.475 1.965 ;
        RECT  0.000 1.635 0.365 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.185 1.040 2.295 1.470 ;
        RECT  0.735 1.210 2.185 1.305 ;
        RECT  0.625 1.040 0.735 1.470 ;
        RECT  0.215 1.040 0.625 1.150 ;
        RECT  0.105 1.040 0.215 1.470 ;
    END
END NR2XD2

MACRO NR2XD3
    CLASS CORE ;
    FOREIGN NR2XD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.010 3.105 1.120 ;
        RECT  2.425 0.270 2.535 0.690 ;
        RECT  2.050 0.575 2.425 0.690 ;
        RECT  1.905 0.270 2.050 1.120 ;
        RECT  1.750 0.575 1.905 1.120 ;
        RECT  1.495 0.575 1.750 0.690 ;
        RECT  1.385 0.270 1.495 0.690 ;
        RECT  0.975 0.575 1.385 0.690 ;
        RECT  0.865 0.270 0.975 0.690 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2574 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.780 1.580 0.890 ;
        RECT  0.250 0.710 0.750 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2574 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 3.150 0.890 ;
        RECT  2.210 0.780 2.650 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 -0.165 3.400 0.165 ;
        RECT  2.165 -0.165 2.275 0.485 ;
        RECT  1.765 -0.165 2.165 0.165 ;
        RECT  1.635 -0.165 1.765 0.485 ;
        RECT  1.235 -0.165 1.635 0.165 ;
        RECT  1.125 -0.165 1.235 0.485 ;
        RECT  0.000 -0.165 1.125 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.445 1.635 3.400 1.965 ;
        RECT  1.445 1.395 1.545 1.505 ;
        RECT  1.335 1.395 1.445 1.965 ;
        RECT  0.975 1.635 1.335 1.965 ;
        RECT  0.865 1.240 0.975 1.965 ;
        RECT  0.455 1.635 0.865 1.965 ;
        RECT  0.345 1.240 0.455 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.150 1.010 3.105 1.120 ;
        RECT  2.425 0.270 2.535 0.690 ;
        RECT  2.150 0.575 2.425 0.690 ;
        RECT  1.495 0.575 1.650 0.690 ;
        RECT  1.385 0.270 1.495 0.690 ;
        RECT  0.975 0.575 1.385 0.690 ;
        RECT  0.865 0.270 0.975 0.690 ;
        RECT  3.205 1.040 3.315 1.470 ;
        RECT  1.235 1.210 3.205 1.305 ;
        RECT  1.125 1.040 1.235 1.470 ;
        RECT  0.715 1.040 1.125 1.150 ;
        RECT  0.605 1.040 0.715 1.470 ;
        RECT  0.195 1.040 0.605 1.150 ;
        RECT  0.085 1.040 0.195 1.470 ;
    END
END NR2XD3

MACRO NR2XD4
    CLASS CORE ;
    FOREIGN NR2XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.140 4.115 1.250 ;
        RECT  2.915 0.270 3.025 0.690 ;
        RECT  2.650 0.575 2.915 0.690 ;
        RECT  2.550 0.575 2.650 1.250 ;
        RECT  2.395 0.270 2.550 1.250 ;
        RECT  2.350 0.575 2.395 1.250 ;
        RECT  1.985 0.575 2.350 0.690 ;
        RECT  1.875 0.270 1.985 0.690 ;
        RECT  1.465 0.575 1.875 0.690 ;
        RECT  1.355 0.270 1.465 0.690 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.3437 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 2.050 0.890 ;
        RECT  0.250 0.710 0.950 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.710 4.150 0.890 ;
        RECT  2.790 0.780 3.450 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.285 -0.165 4.400 0.165 ;
        RECT  3.175 -0.165 3.285 0.690 ;
        RECT  2.765 -0.165 3.175 0.165 ;
        RECT  2.655 -0.165 2.765 0.485 ;
        RECT  2.245 -0.165 2.655 0.165 ;
        RECT  2.135 -0.165 2.245 0.485 ;
        RECT  1.725 -0.165 2.135 0.165 ;
        RECT  1.615 -0.165 1.725 0.485 ;
        RECT  1.205 -0.165 1.615 0.165 ;
        RECT  1.095 -0.165 1.205 0.690 ;
        RECT  0.000 -0.165 1.095 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 1.635 4.400 1.965 ;
        RECT  1.375 1.240 1.485 1.965 ;
        RECT  0.965 1.635 1.375 1.965 ;
        RECT  0.855 1.240 0.965 1.965 ;
        RECT  0.445 1.635 0.855 1.965 ;
        RECT  0.335 1.240 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 1.140 4.115 1.250 ;
        RECT  2.915 0.270 3.025 0.690 ;
        RECT  2.750 0.575 2.915 0.690 ;
        RECT  1.985 0.575 2.250 0.690 ;
        RECT  1.875 0.270 1.985 0.690 ;
        RECT  1.465 0.575 1.875 0.690 ;
        RECT  1.355 0.270 1.465 0.690 ;
        RECT  4.215 1.040 4.325 1.470 ;
        RECT  1.745 1.360 4.215 1.470 ;
        RECT  1.635 1.040 1.745 1.470 ;
        RECT  1.225 1.040 1.635 1.150 ;
        RECT  1.115 1.040 1.225 1.470 ;
        RECT  0.705 1.040 1.115 1.150 ;
        RECT  0.595 1.040 0.705 1.470 ;
        RECT  0.185 1.040 0.595 1.150 ;
        RECT  0.075 1.040 0.185 1.470 ;
    END
END NR2XD4

MACRO NR2XD8
    CLASS CORE ;
    FOREIGN NR2XD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.4560 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 1.140 8.305 1.250 ;
        RECT  6.065 0.270 6.175 0.690 ;
        RECT  5.655 0.575 6.065 0.690 ;
        RECT  5.545 0.270 5.655 0.690 ;
        RECT  5.135 0.575 5.545 0.690 ;
        RECT  5.025 0.270 5.135 0.690 ;
        RECT  4.850 0.575 5.025 0.690 ;
        RECT  4.615 0.575 4.850 1.250 ;
        RECT  4.550 0.270 4.615 1.250 ;
        RECT  4.505 0.270 4.550 0.690 ;
        RECT  4.455 1.140 4.550 1.250 ;
        RECT  4.095 0.575 4.505 0.690 ;
        RECT  3.985 0.270 4.095 0.690 ;
        RECT  3.575 0.575 3.985 0.690 ;
        RECT  3.465 0.270 3.575 0.690 ;
        RECT  3.055 0.575 3.465 0.690 ;
        RECT  2.945 0.270 3.055 0.690 ;
        RECT  2.535 0.575 2.945 0.690 ;
        RECT  2.425 0.270 2.535 0.690 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.6864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.780 4.200 0.890 ;
        RECT  0.250 0.710 1.950 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.710 8.150 0.890 ;
        RECT  5.080 0.780 6.650 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.435 -0.165 8.600 0.165 ;
        RECT  6.325 -0.165 6.435 0.690 ;
        RECT  5.915 -0.165 6.325 0.165 ;
        RECT  5.805 -0.165 5.915 0.485 ;
        RECT  5.395 -0.165 5.805 0.165 ;
        RECT  5.285 -0.165 5.395 0.485 ;
        RECT  4.875 -0.165 5.285 0.165 ;
        RECT  4.765 -0.165 4.875 0.485 ;
        RECT  4.355 -0.165 4.765 0.165 ;
        RECT  4.245 -0.165 4.355 0.485 ;
        RECT  3.835 -0.165 4.245 0.165 ;
        RECT  3.725 -0.165 3.835 0.485 ;
        RECT  3.315 -0.165 3.725 0.165 ;
        RECT  3.205 -0.165 3.315 0.485 ;
        RECT  2.795 -0.165 3.205 0.165 ;
        RECT  2.685 -0.165 2.795 0.485 ;
        RECT  2.275 -0.165 2.685 0.165 ;
        RECT  2.165 -0.165 2.275 0.690 ;
        RECT  0.000 -0.165 2.165 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.095 1.635 8.600 1.965 ;
        RECT  3.985 1.240 4.095 1.965 ;
        RECT  3.575 1.635 3.985 1.965 ;
        RECT  3.465 1.240 3.575 1.965 ;
        RECT  3.055 1.635 3.465 1.965 ;
        RECT  2.945 1.240 3.055 1.965 ;
        RECT  2.535 1.635 2.945 1.965 ;
        RECT  2.425 1.240 2.535 1.965 ;
        RECT  2.015 1.635 2.425 1.965 ;
        RECT  1.905 1.240 2.015 1.965 ;
        RECT  1.495 1.635 1.905 1.965 ;
        RECT  1.385 1.240 1.495 1.965 ;
        RECT  0.975 1.635 1.385 1.965 ;
        RECT  0.865 1.240 0.975 1.965 ;
        RECT  0.455 1.635 0.865 1.965 ;
        RECT  0.345 1.240 0.455 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.950 1.140 8.305 1.250 ;
        RECT  6.065 0.270 6.175 0.690 ;
        RECT  5.655 0.575 6.065 0.690 ;
        RECT  5.545 0.270 5.655 0.690 ;
        RECT  5.135 0.575 5.545 0.690 ;
        RECT  5.025 0.270 5.135 0.690 ;
        RECT  4.950 0.575 5.025 0.690 ;
        RECT  4.095 0.575 4.450 0.690 ;
        RECT  3.985 0.270 4.095 0.690 ;
        RECT  3.575 0.575 3.985 0.690 ;
        RECT  3.465 0.270 3.575 0.690 ;
        RECT  3.055 0.575 3.465 0.690 ;
        RECT  2.945 0.270 3.055 0.690 ;
        RECT  2.535 0.575 2.945 0.690 ;
        RECT  2.425 0.270 2.535 0.690 ;
        RECT  8.405 1.040 8.515 1.470 ;
        RECT  4.365 1.360 8.405 1.470 ;
        RECT  4.245 1.040 4.365 1.470 ;
        RECT  3.835 1.040 4.245 1.150 ;
        RECT  3.725 1.040 3.835 1.470 ;
        RECT  3.315 1.040 3.725 1.150 ;
        RECT  3.205 1.040 3.315 1.470 ;
        RECT  2.795 1.040 3.205 1.150 ;
        RECT  2.685 1.040 2.795 1.470 ;
        RECT  2.275 1.040 2.685 1.150 ;
        RECT  2.165 1.040 2.275 1.470 ;
        RECT  1.755 1.040 2.165 1.150 ;
        RECT  1.645 1.040 1.755 1.470 ;
        RECT  1.235 1.040 1.645 1.150 ;
        RECT  1.125 1.040 1.235 1.470 ;
        RECT  0.715 1.040 1.125 1.150 ;
        RECT  0.605 1.040 0.715 1.470 ;
        RECT  0.195 1.040 0.605 1.150 ;
        RECT  0.085 1.040 0.195 1.470 ;
    END
END NR2XD8

MACRO NR3D0
    CLASS CORE ;
    FOREIGN NR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2050 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.160 ;
        RECT  0.965 0.510 1.050 0.600 ;
        RECT  1.000 1.050 1.050 1.160 ;
        RECT  0.850 1.050 1.000 1.515 ;
        RECT  0.855 0.275 0.965 0.600 ;
        RECT  0.445 0.510 0.855 0.600 ;
        RECT  0.335 0.275 0.445 0.600 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.555 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.800 0.940 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.755 -0.165 1.200 0.165 ;
        RECT  0.645 -0.165 0.755 0.420 ;
        RECT  0.185 -0.165 0.645 0.165 ;
        RECT  0.545 0.310 0.645 0.420 ;
        RECT  0.075 -0.165 0.185 0.480 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.635 1.200 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END NR3D0

MACRO NR3D1
    CLASS CORE ;
    FOREIGN NR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.385 1.150 0.475 ;
        RECT  0.445 1.385 1.040 1.495 ;
        RECT  0.355 1.200 0.445 1.495 ;
        RECT  0.150 1.200 0.355 1.305 ;
        RECT  0.050 0.385 0.150 1.305 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0862 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.780 1.680 0.890 ;
        RECT  1.450 0.585 1.550 0.890 ;
        RECT  0.365 0.585 1.450 0.675 ;
        RECT  0.250 0.585 0.365 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0862 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.775 1.360 1.290 ;
        RECT  0.750 1.200 1.240 1.290 ;
        RECT  0.650 0.785 0.750 1.290 ;
        RECT  0.475 0.785 0.650 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0862 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.910 1.150 1.090 ;
        RECT  0.850 0.785 0.960 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.875 -0.165 1.800 0.165 ;
        RECT  0.665 -0.165 0.875 0.295 ;
        RECT  0.305 -0.165 0.665 0.165 ;
        RECT  0.095 -0.165 0.305 0.295 ;
        RECT  0.000 -0.165 0.095 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.040 1.725 1.965 ;
        RECT  0.245 1.635 1.615 1.965 ;
        RECT  0.055 1.415 0.245 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
END NR3D1

MACRO NR3D2
    CLASS CORE ;
    FOREIGN NR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.750 0.425 2.965 0.525 ;
        RECT  2.750 1.120 2.855 1.230 ;
        RECT  2.650 0.425 2.750 1.230 ;
        RECT  0.475 0.425 2.650 0.525 ;
        RECT  2.145 1.120 2.650 1.230 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1685 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.640 0.955 0.890 ;
        RECT  0.450 0.640 0.845 0.770 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.640 1.755 0.890 ;
        RECT  1.250 0.640 1.645 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1691 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.640 2.555 0.890 ;
        RECT  2.050 0.640 2.445 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.660 -0.165 3.200 0.165 ;
        RECT  2.490 -0.165 2.660 0.335 ;
        RECT  2.090 -0.165 2.490 0.165 ;
        RECT  1.920 -0.165 2.090 0.335 ;
        RECT  1.520 -0.165 1.920 0.165 ;
        RECT  1.350 -0.165 1.520 0.335 ;
        RECT  0.950 -0.165 1.350 0.165 ;
        RECT  0.780 -0.165 0.950 0.335 ;
        RECT  0.375 -0.165 0.780 0.165 ;
        RECT  0.265 -0.165 0.375 0.520 ;
        RECT  0.000 -0.165 0.265 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.995 1.635 3.200 1.965 ;
        RECT  0.885 1.250 0.995 1.965 ;
        RECT  0.475 1.635 0.885 1.965 ;
        RECT  0.365 1.250 0.475 1.965 ;
        RECT  0.000 1.635 0.365 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.965 1.115 3.075 1.460 ;
        RECT  2.035 1.350 2.965 1.460 ;
        RECT  1.925 1.000 2.035 1.460 ;
        RECT  1.355 1.350 1.925 1.460 ;
        RECT  1.255 1.000 1.825 1.110 ;
        RECT  1.145 1.000 1.255 1.460 ;
        RECT  0.735 1.000 1.145 1.110 ;
        RECT  0.625 1.000 0.735 1.430 ;
        RECT  0.215 1.000 0.625 1.110 ;
        RECT  0.105 1.000 0.215 1.430 ;
    END
END NR3D2

MACRO NR3D3
    CLASS CORE ;
    FOREIGN NR3D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7010 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 1.110 4.515 1.240 ;
        RECT  3.650 0.425 4.425 0.525 ;
        RECT  3.350 0.425 3.650 1.240 ;
        RECT  0.250 0.425 3.350 0.525 ;
        RECT  3.265 1.110 3.350 1.240 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.2597 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.620 1.555 0.890 ;
        RECT  0.590 0.620 1.445 0.770 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2597 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.620 2.955 0.890 ;
        RECT  1.990 0.620 2.845 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2598 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.620 4.355 0.890 ;
        RECT  3.850 0.620 4.245 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.645 -0.165 4.800 0.165 ;
        RECT  4.535 -0.165 4.645 0.520 ;
        RECT  4.130 -0.165 4.535 0.165 ;
        RECT  3.960 -0.165 4.130 0.335 ;
        RECT  3.560 -0.165 3.960 0.165 ;
        RECT  3.390 -0.165 3.560 0.335 ;
        RECT  2.990 -0.165 3.390 0.165 ;
        RECT  2.820 -0.165 2.990 0.335 ;
        RECT  2.420 -0.165 2.820 0.165 ;
        RECT  2.250 -0.165 2.420 0.335 ;
        RECT  1.850 -0.165 2.250 0.165 ;
        RECT  1.680 -0.165 1.850 0.335 ;
        RECT  1.280 -0.165 1.680 0.165 ;
        RECT  1.110 -0.165 1.280 0.335 ;
        RECT  0.710 -0.165 1.110 0.165 ;
        RECT  0.540 -0.165 0.710 0.335 ;
        RECT  0.000 -0.165 0.540 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.605 1.635 4.800 1.965 ;
        RECT  1.495 1.250 1.605 1.965 ;
        RECT  1.085 1.635 1.495 1.965 ;
        RECT  0.975 1.250 1.085 1.965 ;
        RECT  0.565 1.635 0.975 1.965 ;
        RECT  0.455 1.000 0.565 1.965 ;
        RECT  0.000 1.635 0.455 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 1.110 4.515 1.240 ;
        RECT  3.750 0.425 4.425 0.525 ;
        RECT  0.250 0.425 3.250 0.525 ;
        RECT  4.615 1.090 4.725 1.460 ;
        RECT  3.165 1.350 4.615 1.460 ;
        RECT  3.055 1.000 3.165 1.460 ;
        RECT  1.965 1.350 3.055 1.460 ;
        RECT  1.865 1.000 2.955 1.110 ;
        RECT  1.755 1.000 1.865 1.460 ;
        RECT  1.345 1.000 1.755 1.110 ;
        RECT  1.235 1.000 1.345 1.460 ;
        RECT  0.825 1.000 1.235 1.110 ;
        RECT  0.715 1.000 0.825 1.460 ;
    END
END NR3D3

MACRO NR3D4
    CLASS CORE ;
    FOREIGN NR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8930 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.615 1.040 5.725 1.480 ;
        RECT  4.650 1.040 5.615 1.230 ;
        RECT  4.650 0.425 5.245 0.525 ;
        RECT  4.350 0.425 4.650 1.230 ;
        RECT  0.475 0.425 4.350 0.525 ;
        RECT  4.005 1.040 4.350 1.230 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.3369 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.620 1.555 0.890 ;
        RECT  0.595 0.620 1.445 0.770 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3373 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.620 3.355 0.890 ;
        RECT  2.395 0.620 3.245 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3375 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.445 0.620 5.555 0.890 ;
        RECT  4.845 0.620 5.445 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.465 -0.165 5.800 0.165 ;
        RECT  5.355 -0.165 5.465 0.520 ;
        RECT  4.950 -0.165 5.355 0.165 ;
        RECT  4.780 -0.165 4.950 0.335 ;
        RECT  4.380 -0.165 4.780 0.165 ;
        RECT  4.210 -0.165 4.380 0.335 ;
        RECT  3.810 -0.165 4.210 0.165 ;
        RECT  3.630 -0.165 3.810 0.335 ;
        RECT  3.230 -0.165 3.630 0.165 ;
        RECT  3.060 -0.165 3.230 0.335 ;
        RECT  2.660 -0.165 3.060 0.165 ;
        RECT  2.490 -0.165 2.660 0.335 ;
        RECT  2.090 -0.165 2.490 0.165 ;
        RECT  1.920 -0.165 2.090 0.335 ;
        RECT  1.520 -0.165 1.920 0.165 ;
        RECT  1.350 -0.165 1.520 0.335 ;
        RECT  0.950 -0.165 1.350 0.165 ;
        RECT  0.780 -0.165 0.950 0.335 ;
        RECT  0.375 -0.165 0.780 0.165 ;
        RECT  0.265 -0.165 0.375 0.520 ;
        RECT  0.000 -0.165 0.265 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.825 1.635 5.800 1.965 ;
        RECT  1.715 1.250 1.825 1.965 ;
        RECT  1.305 1.635 1.715 1.965 ;
        RECT  1.195 1.250 1.305 1.965 ;
        RECT  0.785 1.635 1.195 1.965 ;
        RECT  0.675 1.250 0.785 1.965 ;
        RECT  0.000 1.635 0.675 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.615 1.040 5.725 1.480 ;
        RECT  4.750 1.040 5.615 1.230 ;
        RECT  4.750 0.425 5.245 0.525 ;
        RECT  0.475 0.425 4.250 0.525 ;
        RECT  4.005 1.040 4.250 1.230 ;
        RECT  3.905 1.350 5.515 1.460 ;
        RECT  3.795 1.000 3.905 1.460 ;
        RECT  2.185 1.350 3.795 1.460 ;
        RECT  2.085 1.000 3.675 1.110 ;
        RECT  1.975 1.000 2.085 1.460 ;
        RECT  1.565 1.000 1.975 1.110 ;
        RECT  1.455 1.000 1.565 1.460 ;
        RECT  1.045 1.000 1.455 1.110 ;
        RECT  0.935 1.000 1.045 1.460 ;
        RECT  0.525 1.000 0.935 1.110 ;
        RECT  0.415 1.000 0.525 1.460 ;
    END
END NR3D4

MACRO NR3D8
    CLASS CORE ;
    FOREIGN NR3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.7630 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.215 1.040 10.325 1.480 ;
        RECT  7.650 1.040 10.215 1.230 ;
        RECT  7.650 0.425 10.115 0.525 ;
        RECT  7.350 0.425 7.650 1.230 ;
        RECT  0.285 0.425 7.350 0.525 ;
        RECT  7.045 1.040 7.350 1.230 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.6745 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.620 2.355 0.890 ;
        RECT  1.395 0.620 2.245 0.770 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.6746 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.445 0.620 5.555 0.890 ;
        RECT  4.595 0.620 5.445 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6748 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.045 0.620 9.155 0.890 ;
        RECT  8.195 0.620 9.045 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.325 -0.165 10.400 0.165 ;
        RECT  10.215 -0.165 10.325 0.520 ;
        RECT  9.310 -0.165 10.215 0.165 ;
        RECT  9.140 -0.165 9.310 0.335 ;
        RECT  8.740 -0.165 9.140 0.165 ;
        RECT  8.570 -0.165 8.740 0.335 ;
        RECT  8.170 -0.165 8.570 0.165 ;
        RECT  8.000 -0.165 8.170 0.335 ;
        RECT  7.600 -0.165 8.000 0.165 ;
        RECT  7.430 -0.165 7.600 0.335 ;
        RECT  7.030 -0.165 7.430 0.165 ;
        RECT  6.860 -0.165 7.030 0.335 ;
        RECT  6.460 -0.165 6.860 0.165 ;
        RECT  6.290 -0.165 6.460 0.335 ;
        RECT  5.890 -0.165 6.290 0.165 ;
        RECT  5.720 -0.165 5.890 0.335 ;
        RECT  5.320 -0.165 5.720 0.165 ;
        RECT  5.150 -0.165 5.320 0.335 ;
        RECT  4.750 -0.165 5.150 0.165 ;
        RECT  4.580 -0.165 4.750 0.335 ;
        RECT  4.180 -0.165 4.580 0.165 ;
        RECT  4.010 -0.165 4.180 0.335 ;
        RECT  3.610 -0.165 4.010 0.165 ;
        RECT  3.440 -0.165 3.610 0.335 ;
        RECT  3.040 -0.165 3.440 0.165 ;
        RECT  2.870 -0.165 3.040 0.335 ;
        RECT  2.470 -0.165 2.870 0.165 ;
        RECT  2.300 -0.165 2.470 0.335 ;
        RECT  1.900 -0.165 2.300 0.165 ;
        RECT  1.730 -0.165 1.900 0.335 ;
        RECT  1.330 -0.165 1.730 0.165 ;
        RECT  1.160 -0.165 1.330 0.335 ;
        RECT  0.760 -0.165 1.160 0.165 ;
        RECT  0.590 -0.165 0.760 0.335 ;
        RECT  0.185 -0.165 0.590 0.165 ;
        RECT  0.075 -0.165 0.185 0.520 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 1.635 10.400 1.965 ;
        RECT  3.195 1.250 3.305 1.965 ;
        RECT  2.785 1.635 3.195 1.965 ;
        RECT  2.675 1.250 2.785 1.965 ;
        RECT  2.265 1.635 2.675 1.965 ;
        RECT  2.155 1.250 2.265 1.965 ;
        RECT  1.745 1.635 2.155 1.965 ;
        RECT  1.635 1.250 1.745 1.965 ;
        RECT  1.225 1.635 1.635 1.965 ;
        RECT  1.115 1.250 1.225 1.965 ;
        RECT  0.705 1.635 1.115 1.965 ;
        RECT  0.595 1.250 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.220 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.215 1.040 10.325 1.480 ;
        RECT  7.750 1.040 10.215 1.230 ;
        RECT  7.750 0.425 10.115 0.525 ;
        RECT  0.285 0.425 7.250 0.525 ;
        RECT  7.045 1.040 7.250 1.230 ;
        RECT  6.940 1.350 10.115 1.460 ;
        RECT  6.835 1.000 6.940 1.460 ;
        RECT  3.665 1.350 6.835 1.460 ;
        RECT  3.565 1.000 6.735 1.110 ;
        RECT  3.455 1.000 3.565 1.460 ;
        RECT  3.045 1.000 3.455 1.110 ;
        RECT  2.935 1.000 3.045 1.460 ;
        RECT  2.525 1.000 2.935 1.110 ;
        RECT  2.415 1.000 2.525 1.460 ;
        RECT  2.005 1.000 2.415 1.110 ;
        RECT  1.895 1.000 2.005 1.460 ;
        RECT  1.485 1.000 1.895 1.110 ;
        RECT  1.375 1.000 1.485 1.460 ;
        RECT  0.965 1.000 1.375 1.110 ;
        RECT  0.855 1.000 0.965 1.460 ;
        RECT  0.445 1.000 0.855 1.110 ;
        RECT  0.335 1.000 0.445 1.430 ;
    END
END NR3D8

MACRO NR4D0
    CLASS CORE ;
    FOREIGN NR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.350 1.310 ;
        RECT  0.965 0.510 1.250 0.600 ;
        RECT  1.065 1.200 1.250 1.310 ;
        RECT  0.850 0.285 0.965 0.600 ;
        RECT  0.450 0.510 0.850 0.600 ;
        RECT  0.335 0.285 0.450 0.600 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.350 0.890 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.555 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.790 0.940 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.160 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 -0.165 1.400 0.165 ;
        RECT  1.165 -0.165 1.275 0.400 ;
        RECT  0.755 -0.165 1.165 0.165 ;
        RECT  1.065 0.290 1.165 0.400 ;
        RECT  0.645 -0.165 0.755 0.420 ;
        RECT  0.185 -0.165 0.645 0.165 ;
        RECT  0.545 0.310 0.645 0.420 ;
        RECT  0.075 -0.165 0.185 0.480 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.635 1.400 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
END NR4D0

MACRO NR4D1
    CLASS CORE ;
    FOREIGN NR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1960 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.510 1.715 0.620 ;
        RECT  0.850 0.510 0.950 1.255 ;
        RECT  0.295 0.510 0.850 0.600 ;
        RECT  0.485 1.145 0.850 1.255 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0754 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.710 1.560 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0764 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 0.710 1.950 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0764 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0754 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.925 -0.165 2.000 0.165 ;
        RECT  1.815 -0.165 1.925 0.595 ;
        RECT  1.360 -0.165 1.815 0.165 ;
        RECT  1.190 -0.165 1.360 0.420 ;
        RECT  0.820 -0.165 1.190 0.165 ;
        RECT  0.650 -0.165 0.820 0.420 ;
        RECT  0.195 -0.165 0.650 0.165 ;
        RECT  0.085 -0.165 0.195 0.595 ;
        RECT  0.000 -0.165 0.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.510 1.635 2.000 1.965 ;
        RECT  1.330 1.380 1.510 1.965 ;
        RECT  0.000 1.635 1.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.815 1.200 1.925 1.410 ;
        RECT  1.170 1.200 1.815 1.290 ;
        RECT  1.060 1.200 1.170 1.475 ;
        RECT  0.195 1.365 1.060 1.475 ;
        RECT  0.085 1.265 0.195 1.475 ;
    END
END NR4D1

MACRO NR4D2
    CLASS CORE ;
    FOREIGN NR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5230 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.555 1.120 3.705 1.230 ;
        RECT  3.555 0.425 3.585 0.525 ;
        RECT  3.445 0.425 3.555 1.230 ;
        RECT  0.535 0.425 3.445 0.525 ;
        RECT  2.995 1.120 3.445 1.230 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.1682 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.620 0.950 0.890 ;
        RECT  0.495 0.620 0.850 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.620 1.750 0.890 ;
        RECT  1.250 0.620 1.650 0.770 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.620 2.750 0.890 ;
        RECT  2.250 0.620 2.650 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1687 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.635 3.350 0.890 ;
        RECT  2.955 0.635 3.250 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.795 -0.165 4.000 0.165 ;
        RECT  3.685 -0.165 3.795 0.500 ;
        RECT  3.280 -0.165 3.685 0.165 ;
        RECT  3.110 -0.165 3.280 0.335 ;
        RECT  2.710 -0.165 3.110 0.165 ;
        RECT  2.540 -0.165 2.710 0.335 ;
        RECT  2.140 -0.165 2.540 0.165 ;
        RECT  1.970 -0.165 2.140 0.335 ;
        RECT  1.570 -0.165 1.970 0.165 ;
        RECT  1.400 -0.165 1.570 0.335 ;
        RECT  1.000 -0.165 1.400 0.165 ;
        RECT  0.830 -0.165 1.000 0.335 ;
        RECT  0.425 -0.165 0.830 0.165 ;
        RECT  0.315 -0.165 0.425 0.520 ;
        RECT  0.000 -0.165 0.315 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.065 1.635 4.000 1.965 ;
        RECT  0.955 1.250 1.065 1.965 ;
        RECT  0.545 1.635 0.955 1.965 ;
        RECT  0.435 1.000 0.545 1.965 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.815 1.110 3.925 1.460 ;
        RECT  2.885 1.350 3.815 1.460 ;
        RECT  2.775 1.000 2.885 1.460 ;
        RECT  2.205 1.000 2.775 1.110 ;
        RECT  2.105 1.350 2.675 1.460 ;
        RECT  1.995 1.000 2.105 1.460 ;
        RECT  1.425 1.350 1.995 1.460 ;
        RECT  1.325 1.000 1.895 1.110 ;
        RECT  1.215 1.000 1.325 1.460 ;
        RECT  0.805 1.000 1.215 1.110 ;
        RECT  0.695 1.000 0.805 1.460 ;
    END
END NR4D2

MACRO NR4D3
    CLASS CORE ;
    FOREIGN NR4D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8350 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.805 0.315 5.915 0.525 ;
        RECT  4.850 0.425 5.805 0.525 ;
        RECT  4.850 1.100 5.715 1.210 ;
        RECT  4.550 0.425 4.850 1.210 ;
        RECT  0.055 0.425 4.550 0.525 ;
        RECT  4.465 1.100 4.550 1.210 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.2606 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.620 1.150 0.890 ;
        RECT  0.850 0.710 1.040 0.890 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2597 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 0.620 2.350 0.890 ;
        RECT  2.050 0.710 2.240 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2603 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.840 0.620 3.950 0.890 ;
        RECT  3.650 0.710 3.840 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2632 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.240 0.620 5.350 0.890 ;
        RECT  5.050 0.710 5.240 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 -0.165 6.000 0.165 ;
        RECT  5.490 -0.165 5.660 0.335 ;
        RECT  5.090 -0.165 5.490 0.165 ;
        RECT  4.920 -0.165 5.090 0.335 ;
        RECT  4.510 -0.165 4.920 0.165 ;
        RECT  4.340 -0.165 4.510 0.335 ;
        RECT  3.380 -0.165 4.340 0.165 ;
        RECT  3.210 -0.165 3.380 0.335 ;
        RECT  2.810 -0.165 3.210 0.165 ;
        RECT  2.640 -0.165 2.810 0.335 ;
        RECT  1.710 -0.165 2.640 0.165 ;
        RECT  1.500 -0.165 1.710 0.335 ;
        RECT  1.100 -0.165 1.500 0.165 ;
        RECT  0.930 -0.165 1.100 0.335 ;
        RECT  0.530 -0.165 0.930 0.165 ;
        RECT  0.360 -0.165 0.530 0.335 ;
        RECT  0.000 -0.165 0.360 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 1.635 6.000 1.965 ;
        RECT  1.395 1.220 1.505 1.965 ;
        RECT  0.985 1.635 1.395 1.965 ;
        RECT  0.875 1.220 0.985 1.965 ;
        RECT  0.465 1.635 0.875 1.965 ;
        RECT  0.355 1.220 0.465 1.965 ;
        RECT  0.000 1.635 0.355 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.805 0.315 5.915 0.525 ;
        RECT  4.950 0.425 5.805 0.525 ;
        RECT  4.950 1.100 5.715 1.210 ;
        RECT  0.055 0.425 4.450 0.525 ;
        RECT  5.815 1.095 5.925 1.430 ;
        RECT  4.365 1.320 5.815 1.430 ;
        RECT  4.255 1.000 4.365 1.430 ;
        RECT  3.165 1.000 4.255 1.110 ;
        RECT  3.065 1.320 4.155 1.430 ;
        RECT  2.955 1.000 3.065 1.430 ;
        RECT  1.865 1.320 2.955 1.430 ;
        RECT  1.765 1.000 2.855 1.110 ;
        RECT  1.655 1.000 1.765 1.430 ;
        RECT  1.245 1.000 1.655 1.110 ;
        RECT  1.135 1.000 1.245 1.430 ;
        RECT  0.725 1.000 1.135 1.110 ;
        RECT  0.615 1.000 0.725 1.430 ;
        RECT  0.205 1.000 0.615 1.110 ;
        RECT  0.095 1.000 0.205 1.430 ;
    END
END NR4D3

MACRO NR4D4
    CLASS CORE ;
    FOREIGN NR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.0490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.215 1.040 7.325 1.525 ;
        RECT  6.250 1.040 7.215 1.230 ;
        RECT  6.250 0.425 6.995 0.525 ;
        RECT  5.950 0.425 6.250 1.230 ;
        RECT  0.525 0.425 5.950 0.525 ;
        RECT  5.605 1.040 5.950 1.230 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.3369 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.620 1.555 0.890 ;
        RECT  0.595 0.620 1.445 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.3373 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.620 3.355 0.890 ;
        RECT  2.395 0.620 3.245 0.770 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3373 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.045 0.620 5.155 0.890 ;
        RECT  4.195 0.620 5.045 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3374 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.045 0.620 7.155 0.890 ;
        RECT  6.445 0.620 7.045 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.215 -0.165 7.400 0.165 ;
        RECT  7.105 -0.165 7.215 0.520 ;
        RECT  6.700 -0.165 7.105 0.165 ;
        RECT  6.530 -0.165 6.700 0.335 ;
        RECT  6.130 -0.165 6.530 0.165 ;
        RECT  5.960 -0.165 6.130 0.335 ;
        RECT  5.560 -0.165 5.960 0.165 ;
        RECT  5.390 -0.165 5.560 0.335 ;
        RECT  4.990 -0.165 5.390 0.165 ;
        RECT  4.820 -0.165 4.990 0.335 ;
        RECT  4.420 -0.165 4.820 0.165 ;
        RECT  4.250 -0.165 4.420 0.335 ;
        RECT  3.850 -0.165 4.250 0.165 ;
        RECT  3.670 -0.165 3.850 0.335 ;
        RECT  3.270 -0.165 3.670 0.165 ;
        RECT  3.100 -0.165 3.270 0.335 ;
        RECT  2.700 -0.165 3.100 0.165 ;
        RECT  2.530 -0.165 2.700 0.335 ;
        RECT  2.130 -0.165 2.530 0.165 ;
        RECT  1.960 -0.165 2.130 0.335 ;
        RECT  1.560 -0.165 1.960 0.165 ;
        RECT  1.390 -0.165 1.560 0.335 ;
        RECT  0.990 -0.165 1.390 0.165 ;
        RECT  0.820 -0.165 0.990 0.335 ;
        RECT  0.415 -0.165 0.820 0.165 ;
        RECT  0.305 -0.165 0.415 0.520 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.865 1.635 7.400 1.965 ;
        RECT  1.755 1.250 1.865 1.965 ;
        RECT  1.345 1.635 1.755 1.965 ;
        RECT  1.235 1.250 1.345 1.965 ;
        RECT  0.825 1.635 1.235 1.965 ;
        RECT  0.715 1.250 0.825 1.965 ;
        RECT  0.000 1.635 0.715 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.215 1.040 7.325 1.525 ;
        RECT  6.350 1.040 7.215 1.230 ;
        RECT  6.350 0.425 6.995 0.525 ;
        RECT  0.525 0.425 5.850 0.525 ;
        RECT  5.605 1.040 5.850 1.230 ;
        RECT  3.805 1.370 7.115 1.480 ;
        RECT  2.225 1.000 5.295 1.110 ;
        RECT  2.125 1.350 3.715 1.460 ;
        RECT  2.015 1.000 2.125 1.460 ;
        RECT  1.605 1.000 2.015 1.110 ;
        RECT  1.495 1.000 1.605 1.460 ;
        RECT  1.085 1.000 1.495 1.110 ;
        RECT  0.975 1.000 1.085 1.460 ;
        RECT  0.565 1.000 0.975 1.110 ;
        RECT  0.455 1.000 0.565 1.460 ;
    END
END NR4D4

MACRO NR4D8
    CLASS CORE ;
    FOREIGN NR4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 3.105 0.680 ;
        RECT  2.250 1.015 3.105 1.115 ;
        RECT  1.950 0.510 2.250 1.115 ;
        RECT  1.335 0.510 1.950 0.680 ;
        RECT  1.355 1.015 1.950 1.115 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.165 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.780 0.710 0.850 0.930 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.565 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.835 -0.165 4.200 0.165 ;
        RECT  3.725 -0.165 3.835 0.495 ;
        RECT  3.315 -0.165 3.725 0.165 ;
        RECT  3.205 -0.165 3.315 0.495 ;
        RECT  2.570 -0.165 3.205 0.165 ;
        RECT  2.570 0.305 2.845 0.415 ;
        RECT  2.430 -0.165 2.570 0.415 ;
        RECT  1.570 -0.165 2.430 0.165 ;
        RECT  2.115 0.305 2.430 0.415 ;
        RECT  1.570 0.305 1.805 0.415 ;
        RECT  1.430 -0.165 1.570 0.415 ;
        RECT  0.570 -0.165 1.430 0.165 ;
        RECT  1.075 0.305 1.430 0.415 ;
        RECT  0.570 0.305 0.765 0.415 ;
        RECT  0.430 -0.165 0.570 0.415 ;
        RECT  0.000 -0.165 0.430 0.165 ;
        RECT  0.055 0.305 0.430 0.415 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.635 4.200 1.965 ;
        RECT  3.570 1.385 3.885 1.495 ;
        RECT  3.430 1.385 3.570 1.965 ;
        RECT  3.155 1.385 3.430 1.495 ;
        RECT  2.570 1.635 3.430 1.965 ;
        RECT  2.570 1.385 2.845 1.495 ;
        RECT  2.430 1.385 2.570 1.965 ;
        RECT  2.115 1.385 2.430 1.495 ;
        RECT  1.570 1.635 2.430 1.965 ;
        RECT  1.570 1.385 1.805 1.495 ;
        RECT  1.430 1.385 1.570 1.965 ;
        RECT  1.075 1.385 1.430 1.495 ;
        RECT  0.000 1.635 1.430 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.510 3.105 0.680 ;
        RECT  2.350 1.015 3.105 1.115 ;
        RECT  1.335 0.510 1.850 0.680 ;
        RECT  1.355 1.015 1.850 1.115 ;
        RECT  3.985 0.375 4.095 1.470 ;
        RECT  3.575 0.605 3.985 0.695 ;
        RECT  3.415 1.160 3.985 1.270 ;
        RECT  3.530 0.785 3.870 0.890 ;
        RECT  3.465 0.375 3.575 0.695 ;
        RECT  3.440 0.785 3.530 1.070 ;
        RECT  3.305 0.605 3.465 0.695 ;
        RECT  3.305 0.980 3.440 1.070 ;
        RECT  3.215 0.605 3.305 0.890 ;
        RECT  3.215 0.980 3.305 1.295 ;
        RECT  2.570 0.775 3.215 0.890 ;
        RECT  0.360 1.205 3.215 1.295 ;
        RECT  0.360 0.510 1.025 0.600 ;
        RECT  0.270 0.510 0.360 1.295 ;
        RECT  0.195 1.205 0.270 1.295 ;
        RECT  0.085 1.205 0.195 1.415 ;
    END
END NR4D8

MACRO OA211D0
    CLASS CORE ;
    FOREIGN OA211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.295 1.550 1.495 ;
        RECT  1.375 0.295 1.450 0.405 ;
        RECT  1.375 1.390 1.450 1.495 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.940 0.780 1.050 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.840 0.940 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 -0.165 1.600 0.165 ;
        RECT  1.175 -0.165 1.285 0.405 ;
        RECT  0.000 -0.165 1.175 0.165 ;
        RECT  1.095 0.295 1.175 0.405 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.175 1.635 1.600 1.965 ;
        RECT  1.175 1.390 1.265 1.500 ;
        RECT  1.065 1.390 1.175 1.965 ;
        RECT  0.755 1.635 1.065 1.965 ;
        RECT  0.645 1.390 0.755 1.965 ;
        RECT  0.545 1.390 0.645 1.500 ;
        RECT  0.000 1.635 0.645 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.495 1.340 1.300 ;
        RECT  0.310 0.495 1.240 0.600 ;
        RECT  0.965 1.200 1.240 1.300 ;
        RECT  0.855 1.200 0.965 1.490 ;
        RECT  0.185 1.200 0.855 1.300 ;
        RECT  0.175 0.295 0.805 0.405 ;
        RECT  0.075 1.200 0.185 1.490 ;
        RECT  0.075 0.295 0.175 0.505 ;
    END
END OA211D0

MACRO OA211D1
    CLASS CORE ;
    FOREIGN OA211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.305 1.550 1.495 ;
        RECT  1.365 0.305 1.450 0.410 ;
        RECT  1.365 1.390 1.450 1.495 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.900 0.780 1.050 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.790 0.940 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.255 -0.165 1.600 0.165 ;
        RECT  1.085 -0.165 1.255 0.410 ;
        RECT  0.000 -0.165 1.085 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.635 1.600 1.965 ;
        RECT  0.970 1.390 1.255 1.495 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.545 1.390 0.830 1.495 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.500 1.340 1.300 ;
        RECT  0.285 0.500 1.240 0.600 ;
        RECT  0.185 1.200 1.240 1.300 ;
        RECT  0.175 0.305 0.755 0.410 ;
        RECT  0.075 1.200 0.185 1.410 ;
        RECT  0.075 0.305 0.175 0.520 ;
    END
END OA211D1

MACRO OA211D2
    CLASS CORE ;
    FOREIGN OA211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.290 ;
        RECT  1.315 0.510 1.450 0.620 ;
        RECT  1.305 1.180 1.450 1.290 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.890 ;
        RECT  0.940 0.780 1.050 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.800 0.940 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.560 1.095 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.445 ;
        RECT  1.205 -0.165 1.615 0.165 ;
        RECT  1.035 -0.165 1.205 0.410 ;
        RECT  0.000 -0.165 1.035 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.355 1.725 1.965 ;
        RECT  0.970 1.635 1.615 1.965 ;
        RECT  0.970 1.390 1.255 1.495 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.525 1.390 0.830 1.495 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.755 1.340 1.090 ;
        RECT  1.195 1.000 1.240 1.090 ;
        RECT  1.105 1.000 1.195 1.300 ;
        RECT  0.360 1.205 1.105 1.300 ;
        RECT  0.175 0.300 0.755 0.400 ;
        RECT  0.360 0.510 0.495 0.600 ;
        RECT  0.270 0.510 0.360 1.300 ;
        RECT  0.185 1.200 0.270 1.300 ;
        RECT  0.075 1.200 0.185 1.410 ;
        RECT  0.075 0.300 0.175 0.520 ;
    END
END OA211D2

MACRO OA211D4
    CLASS CORE ;
    FOREIGN OA211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.155 0.275 3.265 0.675 ;
        RECT  3.155 1.040 3.265 1.470 ;
        RECT  3.050 0.585 3.155 0.675 ;
        RECT  3.050 1.040 3.155 1.150 ;
        RECT  2.750 0.585 3.050 1.150 ;
        RECT  2.635 0.275 2.750 0.675 ;
        RECT  2.635 1.040 2.750 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.710 1.150 0.890 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.180 1.000 0.850 1.090 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.710 2.060 1.090 ;
        RECT  1.350 1.000 1.950 1.090 ;
        RECT  1.250 0.710 1.350 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 -0.165 3.600 0.165 ;
        RECT  3.415 -0.165 3.525 0.695 ;
        RECT  3.005 -0.165 3.415 0.165 ;
        RECT  2.895 -0.165 3.005 0.475 ;
        RECT  2.485 -0.165 2.895 0.165 ;
        RECT  2.375 -0.165 2.485 0.675 ;
        RECT  0.740 -0.165 2.375 0.165 ;
        RECT  0.560 -0.165 0.740 0.420 ;
        RECT  0.000 -0.165 0.560 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 1.635 3.600 1.965 ;
        RECT  3.415 1.040 3.525 1.965 ;
        RECT  3.005 1.635 3.415 1.965 ;
        RECT  2.895 1.260 3.005 1.965 ;
        RECT  2.485 1.635 2.895 1.965 ;
        RECT  2.375 1.040 2.485 1.965 ;
        RECT  2.235 1.635 2.375 1.965 ;
        RECT  2.025 1.415 2.235 1.965 ;
        RECT  0.970 1.635 2.025 1.965 ;
        RECT  0.970 1.390 1.275 1.495 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.545 1.390 0.830 1.495 ;
        RECT  0.185 1.635 0.830 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.155 0.275 3.265 0.675 ;
        RECT  3.155 1.040 3.265 1.470 ;
        RECT  3.150 0.585 3.155 0.675 ;
        RECT  3.150 1.040 3.155 1.150 ;
        RECT  2.635 0.275 2.650 0.675 ;
        RECT  2.635 1.040 2.650 1.490 ;
        RECT  2.260 0.785 2.630 0.890 ;
        RECT  1.185 0.305 2.265 0.410 ;
        RECT  2.170 0.500 2.260 1.300 ;
        RECT  1.295 0.500 2.170 0.600 ;
        RECT  0.295 1.200 2.170 1.300 ;
        RECT  1.075 0.305 1.185 0.600 ;
        RECT  0.065 0.510 1.075 0.600 ;
    END
END OA211D4

MACRO OA21D0
    CLASS CORE ;
    FOREIGN OA21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.275 1.350 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.860 0.970 ;
        RECT  0.650 0.710 0.750 1.120 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.085 -0.165 1.400 0.165 ;
        RECT  0.905 -0.165 1.085 0.410 ;
        RECT  0.000 -0.165 0.905 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.635 1.400 1.965 ;
        RECT  0.880 1.455 1.030 1.965 ;
        RECT  0.195 1.635 0.880 1.965 ;
        RECT  0.085 1.280 0.195 1.965 ;
        RECT  0.000 1.635 0.085 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.500 1.105 1.340 ;
        RECT  0.320 0.500 1.000 0.600 ;
        RECT  0.715 1.240 1.000 1.340 ;
        RECT  0.190 0.300 0.815 0.410 ;
        RECT  0.605 1.240 0.715 1.490 ;
        RECT  0.070 0.300 0.190 0.510 ;
    END
END OA21D0

MACRO OA21D1
    CLASS CORE ;
    FOREIGN OA21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.275 1.350 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.970 ;
        RECT  0.650 0.700 0.750 1.120 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 -0.165 1.400 0.165 ;
        RECT  0.870 -0.165 1.040 0.410 ;
        RECT  0.000 -0.165 0.870 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.635 1.400 1.965 ;
        RECT  0.870 1.430 1.040 1.965 ;
        RECT  0.190 1.635 0.870 1.965 ;
        RECT  0.070 1.325 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.005 0.500 1.105 1.340 ;
        RECT  0.305 0.500 1.005 0.590 ;
        RECT  0.565 1.240 1.005 1.340 ;
        RECT  0.190 0.310 0.755 0.410 ;
        RECT  0.070 0.310 0.190 0.560 ;
    END
END OA21D1

MACRO OA21D2
    CLASS CORE ;
    FOREIGN OA21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.535 1.350 1.195 ;
        RECT  1.250 0.295 1.260 1.475 ;
        RECT  1.160 0.295 1.250 0.675 ;
        RECT  1.160 1.055 1.250 1.475 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.970 ;
        RECT  0.650 0.700 0.750 1.120 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.530 -0.165 1.600 0.165 ;
        RECT  1.410 -0.165 1.530 0.455 ;
        RECT  1.045 -0.165 1.410 0.165 ;
        RECT  0.855 -0.165 1.045 0.410 ;
        RECT  0.000 -0.165 0.855 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.530 1.635 1.600 1.965 ;
        RECT  1.410 1.325 1.530 1.965 ;
        RECT  1.010 1.635 1.410 1.965 ;
        RECT  0.840 1.430 1.010 1.965 ;
        RECT  0.190 1.635 0.840 1.965 ;
        RECT  0.070 1.325 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.500 1.050 1.340 ;
        RECT  0.305 0.500 0.950 0.590 ;
        RECT  0.545 1.240 0.950 1.340 ;
        RECT  0.190 0.310 0.745 0.410 ;
        RECT  0.070 0.310 0.190 0.560 ;
    END
END OA21D2

MACRO OA21D4
    CLASS CORE ;
    FOREIGN OA21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.430 2.885 0.620 ;
        RECT  2.650 1.105 2.885 1.295 ;
        RECT  2.350 0.430 2.650 1.295 ;
        RECT  2.145 0.430 2.350 0.620 ;
        RECT  2.145 1.105 2.350 1.295 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.700 0.360 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.350 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.560 1.100 ;
        RECT  0.950 1.010 1.450 1.100 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.770 0.700 0.850 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 -0.165 3.200 0.165 ;
        RECT  3.010 -0.165 3.130 0.560 ;
        RECT  2.610 -0.165 3.010 0.165 ;
        RECT  2.420 -0.165 2.610 0.320 ;
        RECT  2.010 -0.165 2.420 0.165 ;
        RECT  1.910 -0.165 2.010 0.560 ;
        RECT  0.485 -0.165 1.910 0.165 ;
        RECT  0.295 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.295 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.635 3.200 1.965 ;
        RECT  3.010 1.240 3.130 1.965 ;
        RECT  2.600 1.635 3.010 1.965 ;
        RECT  2.430 1.385 2.600 1.965 ;
        RECT  2.010 1.635 2.430 1.965 ;
        RECT  1.910 1.240 2.010 1.965 ;
        RECT  0.770 1.635 1.910 1.965 ;
        RECT  0.770 1.390 1.265 1.490 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.295 1.390 0.630 1.490 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 0.430 2.885 0.620 ;
        RECT  2.750 1.105 2.885 1.295 ;
        RECT  2.145 0.430 2.250 0.620 ;
        RECT  2.145 1.105 2.250 1.295 ;
        RECT  1.785 0.780 2.240 0.890 ;
        RECT  0.700 0.310 1.785 0.410 ;
        RECT  1.685 0.500 1.785 1.300 ;
        RECT  0.815 0.500 1.685 0.590 ;
        RECT  0.180 1.210 1.685 1.300 ;
        RECT  0.600 0.310 0.700 0.590 ;
        RECT  0.180 0.500 0.600 0.590 ;
        RECT  0.060 0.350 0.180 0.590 ;
        RECT  0.060 1.210 0.180 1.450 ;
    END
END OA21D4

MACRO OA221D0
    CLASS CORE ;
    FOREIGN OA221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.825 0.445 1.950 1.515 ;
        RECT  1.810 1.345 1.825 1.515 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.690 1.550 1.090 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.710 1.350 1.090 ;
        RECT  1.050 0.835 1.245 0.945 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.895 1.095 1.150 1.270 ;
        RECT  0.160 1.180 0.895 1.270 ;
        RECT  0.050 0.565 0.160 1.270 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 0.855 0.835 0.945 ;
        RECT  0.450 0.855 0.780 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.680 0.360 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 2.000 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.720 0.495 1.735 1.255 ;
        RECT  1.640 0.495 1.720 1.490 ;
        RECT  0.710 0.495 1.640 0.600 ;
        RECT  1.620 1.165 1.640 1.490 ;
        RECT  0.255 1.380 1.620 1.490 ;
        RECT  0.210 0.275 1.365 0.385 ;
        RECT  0.580 0.495 0.710 0.720 ;
        RECT  0.080 0.275 0.210 0.455 ;
    END
END OA221D0

MACRO OA221D1
    CLASS CORE ;
    FOREIGN OA221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.275 2.150 1.490 ;
        RECT  2.005 0.275 2.050 0.675 ;
        RECT  2.005 1.265 2.050 1.490 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.500 1.750 0.910 ;
        RECT  1.580 0.740 1.650 0.910 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.700 1.410 0.950 ;
        RECT  1.250 0.700 1.350 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.700 1.150 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.700 0.755 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.860 -0.165 2.200 0.165 ;
        RECT  1.695 -0.165 1.860 0.390 ;
        RECT  0.000 -0.165 1.695 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.635 2.200 1.965 ;
        RECT  1.690 1.410 1.860 1.965 ;
        RECT  1.050 1.635 1.690 1.965 ;
        RECT  0.880 1.410 1.050 1.965 ;
        RECT  0.250 1.635 0.880 1.965 ;
        RECT  0.080 1.410 0.250 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 0.775 1.940 1.120 ;
        RECT  1.745 1.030 1.840 1.120 ;
        RECT  1.655 1.030 1.745 1.300 ;
        RECT  0.360 1.210 1.655 1.300 ;
        RECT  0.875 0.310 1.585 0.410 ;
        RECT  0.740 0.500 1.325 0.590 ;
        RECT  0.640 0.310 0.740 0.590 ;
        RECT  0.075 0.310 0.640 0.410 ;
        RECT  0.360 0.500 0.525 0.590 ;
        RECT  0.260 0.500 0.360 1.300 ;
    END
END OA221D1

MACRO OA221D2
    CLASS CORE ;
    FOREIGN OA221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.535 2.150 1.195 ;
        RECT  2.050 0.275 2.065 1.475 ;
        RECT  1.955 0.275 2.050 0.675 ;
        RECT  1.955 1.045 2.050 1.475 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.630 0.950 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.360 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.700 1.010 0.950 ;
        RECT  0.850 0.700 0.950 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.165 2.400 0.165 ;
        RECT  2.210 -0.165 2.330 0.455 ;
        RECT  1.820 -0.165 2.210 0.165 ;
        RECT  1.685 -0.165 1.820 0.580 ;
        RECT  0.000 -0.165 1.685 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.635 2.400 1.965 ;
        RECT  2.210 1.325 2.330 1.965 ;
        RECT  1.810 1.635 2.210 1.965 ;
        RECT  1.640 1.410 1.810 1.965 ;
        RECT  1.030 1.635 1.640 1.965 ;
        RECT  0.860 1.410 1.030 1.965 ;
        RECT  0.250 1.635 0.860 1.965 ;
        RECT  0.080 1.410 0.250 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.840 0.775 1.910 0.945 ;
        RECT  1.740 0.775 1.840 1.300 ;
        RECT  0.360 1.210 1.740 1.300 ;
        RECT  0.875 0.310 1.595 0.410 ;
        RECT  0.740 0.500 1.325 0.590 ;
        RECT  0.640 0.310 0.740 0.590 ;
        RECT  0.075 0.310 0.640 0.410 ;
        RECT  0.360 0.500 0.525 0.590 ;
        RECT  0.260 0.500 0.360 1.300 ;
    END
END OA221D2

MACRO OA221D4
    CLASS CORE ;
    FOREIGN OA221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.430 4.105 0.620 ;
        RECT  4.050 1.105 4.105 1.295 ;
        RECT  3.750 0.430 4.050 1.295 ;
        RECT  3.435 0.430 3.750 0.620 ;
        RECT  3.435 1.105 3.750 1.295 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  0.950 1.000 1.650 1.090 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.765 0.710 0.850 0.920 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.750 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.950 1.090 ;
        RECT  2.150 1.000 2.850 1.090 ;
        RECT  2.040 0.710 2.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.165 4.400 0.165 ;
        RECT  4.215 -0.165 4.325 0.695 ;
        RECT  0.485 -0.165 4.215 0.165 ;
        RECT  0.305 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.040 4.325 1.965 ;
        RECT  2.605 1.635 4.215 1.965 ;
        RECT  2.425 1.390 2.605 1.965 ;
        RECT  0.970 1.635 2.425 1.965 ;
        RECT  0.970 1.390 1.280 1.500 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.300 1.390 0.830 1.500 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.435 0.430 3.650 0.620 ;
        RECT  3.435 1.105 3.650 1.295 ;
        RECT  3.185 0.780 3.560 0.890 ;
        RECT  3.085 0.500 3.185 1.300 ;
        RECT  1.900 0.500 3.085 0.600 ;
        RECT  0.190 1.200 3.085 1.300 ;
        RECT  0.810 0.310 2.880 0.410 ;
        RECT  0.190 0.500 1.790 0.600 ;
        RECT  0.065 0.350 0.190 0.600 ;
        RECT  0.065 1.200 0.190 1.450 ;
    END
END OA221D4

MACRO OA222D0
    CLASS CORE ;
    FOREIGN OA222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.275 2.350 1.490 ;
        RECT  2.215 0.275 2.250 0.475 ;
        RECT  2.210 1.265 2.250 1.490 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.710 1.555 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.710 1.880 0.950 ;
        RECT  1.650 0.710 1.750 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.080 -0.165 2.400 0.165 ;
        RECT  1.940 -0.165 2.080 0.480 ;
        RECT  0.000 -0.165 1.940 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.100 1.635 2.400 1.965 ;
        RECT  1.920 1.390 2.100 1.965 ;
        RECT  1.270 1.635 1.920 1.965 ;
        RECT  1.095 1.390 1.270 1.965 ;
        RECT  0.230 1.635 1.095 1.965 ;
        RECT  0.060 1.390 0.230 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.100 0.775 2.150 0.945 ;
        RECT  2.000 0.775 2.100 1.300 ;
        RECT  1.555 1.210 2.000 1.300 ;
        RECT  1.695 0.280 1.805 0.600 ;
        RECT  0.885 0.500 1.695 0.600 ;
        RECT  1.425 1.210 1.555 1.490 ;
        RECT  0.730 1.210 1.425 1.300 ;
        RECT  0.050 0.300 1.380 0.410 ;
        RECT  0.600 1.210 0.730 1.490 ;
        RECT  0.350 1.210 0.600 1.300 ;
        RECT  0.350 0.500 0.525 0.600 ;
        RECT  0.260 0.500 0.350 1.300 ;
    END
END OA222D0

MACRO OA222D1
    CLASS CORE ;
    FOREIGN OA222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.275 2.350 1.490 ;
        RECT  2.205 0.275 2.250 0.675 ;
        RECT  2.210 1.045 2.250 1.490 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.700 1.880 0.950 ;
        RECT  1.650 0.700 1.750 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.155 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 -0.165 2.400 0.165 ;
        RECT  1.945 -0.165 2.055 0.585 ;
        RECT  1.570 -0.165 1.945 0.165 ;
        RECT  1.395 -0.165 1.570 0.410 ;
        RECT  0.000 -0.165 1.395 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.060 1.635 2.400 1.965 ;
        RECT  1.890 1.410 2.060 1.965 ;
        RECT  1.280 1.635 1.890 1.965 ;
        RECT  1.095 1.390 1.280 1.965 ;
        RECT  0.235 1.635 1.095 1.965 ;
        RECT  0.060 1.390 0.235 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.100 0.775 2.140 0.945 ;
        RECT  2.000 0.775 2.100 1.300 ;
        RECT  0.350 1.210 2.000 1.300 ;
        RECT  0.830 0.500 1.835 0.590 ;
        RECT  0.060 0.310 1.270 0.410 ;
        RECT  0.350 0.500 0.500 0.590 ;
        RECT  0.260 0.500 0.350 1.300 ;
    END
END OA222D1

MACRO OA222D2
    CLASS CORE ;
    FOREIGN OA222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.265 0.535 2.350 1.195 ;
        RECT  2.260 0.275 2.265 1.195 ;
        RECT  2.250 0.275 2.260 1.465 ;
        RECT  2.155 0.275 2.250 0.675 ;
        RECT  2.160 1.045 2.250 1.465 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.710 1.555 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.710 1.830 0.960 ;
        RECT  1.650 0.710 1.750 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.960 ;
        RECT  0.650 0.710 0.750 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.155 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.560 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.165 2.600 0.165 ;
        RECT  2.410 -0.165 2.530 0.455 ;
        RECT  2.020 -0.165 2.410 0.165 ;
        RECT  1.885 -0.165 2.020 0.590 ;
        RECT  0.000 -0.165 1.885 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 1.635 2.600 1.965 ;
        RECT  2.410 1.325 2.530 1.965 ;
        RECT  2.010 1.635 2.410 1.965 ;
        RECT  1.840 1.410 2.010 1.965 ;
        RECT  1.245 1.635 1.840 1.965 ;
        RECT  1.060 1.390 1.245 1.965 ;
        RECT  0.240 1.635 1.060 1.965 ;
        RECT  0.060 1.390 0.240 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.050 0.775 2.090 0.945 ;
        RECT  1.950 0.775 2.050 1.300 ;
        RECT  0.360 1.210 1.950 1.300 ;
        RECT  0.815 0.510 1.795 0.600 ;
        RECT  0.705 0.310 1.275 0.420 ;
        RECT  0.595 0.310 0.705 0.570 ;
        RECT  0.180 0.310 0.595 0.400 ;
        RECT  0.360 0.510 0.495 0.600 ;
        RECT  0.270 0.510 0.360 1.300 ;
        RECT  0.075 0.310 0.180 0.570 ;
    END
END OA222D2

MACRO OA222D4
    CLASS CORE ;
    FOREIGN OA222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 0.275 4.635 0.695 ;
        RECT  4.520 1.040 4.635 1.470 ;
        RECT  4.450 0.585 4.520 0.695 ;
        RECT  4.450 1.040 4.520 1.150 ;
        RECT  4.150 0.585 4.450 1.150 ;
        RECT  4.115 0.585 4.150 0.695 ;
        RECT  4.115 1.040 4.150 1.150 ;
        RECT  4.005 0.275 4.115 0.695 ;
        RECT  3.985 1.040 4.115 1.470 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.700 1.150 1.100 ;
        RECT  0.170 1.010 1.030 1.100 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.950 0.900 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.700 2.150 1.100 ;
        RECT  1.370 1.010 2.050 1.100 ;
        RECT  1.250 0.700 1.370 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.700 3.150 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.700 3.420 0.920 ;
        RECT  3.250 0.700 3.350 1.100 ;
        RECT  2.550 1.010 3.250 1.100 ;
        RECT  2.450 0.700 2.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.895 -0.165 5.000 0.165 ;
        RECT  4.785 -0.165 4.895 0.695 ;
        RECT  4.375 -0.165 4.785 0.165 ;
        RECT  4.265 -0.165 4.375 0.475 ;
        RECT  3.855 -0.165 4.265 0.165 ;
        RECT  3.750 -0.165 3.855 0.675 ;
        RECT  0.770 -0.165 3.750 0.165 ;
        RECT  0.770 0.305 1.015 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.295 0.305 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.895 1.635 5.000 1.965 ;
        RECT  4.785 1.040 4.895 1.965 ;
        RECT  4.375 1.635 4.785 1.965 ;
        RECT  4.265 1.260 4.375 1.965 ;
        RECT  3.855 1.635 4.265 1.965 ;
        RECT  3.750 1.040 3.855 1.965 ;
        RECT  2.370 1.635 3.750 1.965 ;
        RECT  2.370 1.390 3.125 1.495 ;
        RECT  2.230 1.390 2.370 1.965 ;
        RECT  1.065 1.390 2.230 1.495 ;
        RECT  0.185 1.635 2.230 1.965 ;
        RECT  0.075 1.230 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.550 0.275 4.635 0.695 ;
        RECT  4.550 1.040 4.635 1.470 ;
        RECT  4.005 0.275 4.050 0.695 ;
        RECT  3.985 1.040 4.050 1.470 ;
        RECT  3.640 0.785 4.040 0.890 ;
        RECT  3.550 0.500 3.640 1.300 ;
        RECT  2.415 0.500 3.550 0.590 ;
        RECT  0.555 1.210 3.550 1.300 ;
        RECT  1.325 0.305 3.385 0.410 ;
        RECT  0.185 0.500 2.305 0.590 ;
        RECT  0.075 0.345 0.185 0.590 ;
    END
END OA222D4

MACRO OA22D0
    CLASS CORE ;
    FOREIGN OA22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.285 1.550 1.515 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.160 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.695 1.150 1.300 ;
        RECT  0.550 1.205 1.045 1.300 ;
        RECT  0.420 1.035 0.550 1.300 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.710 0.950 1.115 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.895 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.245 0.495 1.335 1.490 ;
        RECT  0.580 0.495 1.245 0.585 ;
        RECT  0.470 1.390 1.245 1.490 ;
        RECT  0.290 0.305 1.035 0.405 ;
    END
END OA22D0

MACRO OA22D1
    CLASS CORE ;
    FOREIGN OA22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 0.275 1.750 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.930 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.710 1.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 -0.165 1.800 0.165 ;
        RECT  0.410 0.300 0.510 0.410 ;
        RECT  0.300 -0.165 0.410 0.410 ;
        RECT  0.000 -0.165 0.300 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.755 1.635 1.800 1.965 ;
        RECT  0.575 1.390 0.755 1.965 ;
        RECT  0.000 1.635 0.575 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.320 1.490 1.300 ;
        RECT  0.820 0.320 1.390 0.410 ;
        RECT  0.050 1.200 1.390 1.300 ;
        RECT  0.050 0.500 1.280 0.600 ;
    END
END OA22D1

MACRO OA22D2
    CLASS CORE ;
    FOREIGN OA22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 0.535 1.950 1.195 ;
        RECT  1.850 0.285 1.870 1.465 ;
        RECT  1.750 0.285 1.850 0.675 ;
        RECT  1.750 1.035 1.850 1.465 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.550 1.120 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.120 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.970 ;
        RECT  0.650 0.700 0.750 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 -0.165 2.200 0.165 ;
        RECT  2.010 -0.165 2.130 0.455 ;
        RECT  1.610 -0.165 2.010 0.165 ;
        RECT  1.440 -0.165 1.610 0.390 ;
        RECT  0.500 -0.165 1.440 0.165 ;
        RECT  0.310 -0.165 0.500 0.410 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 1.635 2.200 1.965 ;
        RECT  2.010 1.325 2.130 1.965 ;
        RECT  1.610 1.635 2.010 1.965 ;
        RECT  1.440 1.455 1.610 1.965 ;
        RECT  0.750 1.635 1.440 1.965 ;
        RECT  0.580 1.455 0.750 1.965 ;
        RECT  0.000 1.635 0.580 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.500 0.500 1.600 1.340 ;
        RECT  0.830 0.500 1.500 0.590 ;
        RECT  0.060 1.240 1.500 1.340 ;
        RECT  0.715 0.310 1.280 0.410 ;
        RECT  0.615 0.310 0.715 0.590 ;
        RECT  0.195 0.500 0.615 0.590 ;
        RECT  0.075 0.350 0.195 0.590 ;
    END
END OA22D2

MACRO OA22D4
    CLASS CORE ;
    FOREIGN OA22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.275 3.265 0.695 ;
        RECT  3.150 1.040 3.265 1.470 ;
        RECT  3.050 0.585 3.150 0.695 ;
        RECT  3.050 1.040 3.150 1.150 ;
        RECT  2.750 0.585 3.050 1.150 ;
        RECT  2.745 0.585 2.750 0.695 ;
        RECT  2.745 1.040 2.750 1.150 ;
        RECT  2.635 0.275 2.745 0.695 ;
        RECT  2.615 1.040 2.745 1.470 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.710 1.065 1.090 ;
        RECT  0.180 1.000 0.955 1.090 ;
        RECT  0.050 0.700 0.180 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.710 0.750 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.710 2.050 0.940 ;
        RECT  1.850 0.710 1.950 1.090 ;
        RECT  1.350 1.000 1.850 1.090 ;
        RECT  1.225 0.710 1.350 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 -0.165 3.600 0.165 ;
        RECT  3.415 -0.165 3.525 0.695 ;
        RECT  3.005 -0.165 3.415 0.165 ;
        RECT  2.895 -0.165 3.005 0.475 ;
        RECT  2.485 -0.165 2.895 0.165 ;
        RECT  2.375 -0.165 2.485 0.675 ;
        RECT  0.000 -0.165 2.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 1.635 3.600 1.965 ;
        RECT  3.415 1.040 3.525 1.965 ;
        RECT  3.005 1.635 3.415 1.965 ;
        RECT  2.895 1.260 3.005 1.965 ;
        RECT  2.485 1.635 2.895 1.965 ;
        RECT  2.375 1.040 2.485 1.965 ;
        RECT  1.770 1.635 2.375 1.965 ;
        RECT  1.770 1.390 2.265 1.490 ;
        RECT  1.630 1.390 1.770 1.965 ;
        RECT  1.025 1.390 1.630 1.490 ;
        RECT  0.185 1.635 1.630 1.965 ;
        RECT  0.075 1.210 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 0.275 3.265 0.695 ;
        RECT  3.150 1.040 3.265 1.470 ;
        RECT  2.635 0.275 2.650 0.695 ;
        RECT  2.615 1.040 2.650 1.470 ;
        RECT  2.265 0.785 2.640 0.890 ;
        RECT  0.715 0.310 2.265 0.410 ;
        RECT  2.165 0.500 2.265 1.300 ;
        RECT  1.285 0.500 2.165 0.600 ;
        RECT  0.525 1.200 2.165 1.300 ;
        RECT  0.545 0.310 0.715 0.610 ;
        RECT  0.185 0.310 0.545 0.410 ;
        RECT  0.075 0.310 0.185 0.585 ;
    END
END OA22D4

MACRO OA31D0
    CLASS CORE ;
    FOREIGN OA31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.295 1.550 1.490 ;
        RECT  1.405 0.295 1.450 0.485 ;
        RECT  1.405 1.265 1.450 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.500 1.150 0.910 ;
        RECT  1.000 0.740 1.030 0.910 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.790 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.635 1.600 1.965 ;
        RECT  1.090 1.455 1.260 1.965 ;
        RECT  0.235 1.635 1.090 1.965 ;
        RECT  0.055 1.390 0.235 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.730 1.360 1.120 ;
        RECT  1.145 1.030 1.250 1.120 ;
        RECT  1.055 1.030 1.145 1.300 ;
        RECT  0.285 0.300 1.065 0.410 ;
        RECT  0.945 1.210 1.055 1.300 ;
        RECT  0.835 1.210 0.945 1.490 ;
        RECT  0.350 1.210 0.835 1.300 ;
        RECT  0.350 0.500 0.775 0.600 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.075 0.280 0.185 0.590 ;
    END
END OA31D0

MACRO OA31D1
    CLASS CORE ;
    FOREIGN OA31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.295 1.550 1.490 ;
        RECT  1.405 0.295 1.450 0.675 ;
        RECT  1.405 1.265 1.450 1.490 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.500 1.150 0.910 ;
        RECT  0.950 0.740 1.030 0.910 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.700 0.790 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 -0.165 1.600 0.165 ;
        RECT  1.105 -0.165 1.285 0.410 ;
        RECT  0.000 -0.165 1.105 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.635 1.600 1.965 ;
        RECT  1.090 1.455 1.260 1.965 ;
        RECT  0.235 1.635 1.090 1.965 ;
        RECT  0.055 1.390 0.235 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.775 1.340 1.120 ;
        RECT  1.145 1.030 1.240 1.120 ;
        RECT  1.055 1.030 1.145 1.300 ;
        RECT  0.350 1.210 1.055 1.300 ;
        RECT  0.295 0.310 0.995 0.410 ;
        RECT  0.350 0.500 0.745 0.590 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 0.500 0.260 0.590 ;
        RECT  0.060 0.350 0.180 0.590 ;
    END
END OA31D1

MACRO OA31D2
    CLASS CORE ;
    FOREIGN OA31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.465 0.575 1.550 1.300 ;
        RECT  1.450 0.275 1.465 1.300 ;
        RECT  1.355 0.275 1.450 0.665 ;
        RECT  1.305 1.200 1.450 1.300 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.510 1.150 0.890 ;
        RECT  0.900 0.765 1.030 0.890 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.790 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.555 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.465 ;
        RECT  0.000 -0.165 1.615 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 1.635 1.800 1.965 ;
        RECT  1.580 1.390 1.755 1.965 ;
        RECT  1.240 1.635 1.580 1.965 ;
        RECT  1.060 1.390 1.240 1.965 ;
        RECT  0.220 1.635 1.060 1.965 ;
        RECT  0.045 1.390 0.220 1.965 ;
        RECT  0.000 1.635 0.045 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.775 1.360 1.070 ;
        RECT  1.145 0.980 1.260 1.070 ;
        RECT  1.055 0.980 1.145 1.300 ;
        RECT  0.350 1.200 1.055 1.300 ;
        RECT  0.295 0.310 1.015 0.410 ;
        RECT  0.350 0.500 0.755 0.600 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.045 0.500 0.260 0.600 ;
    END
END OA31D2

MACRO OA31D4
    CLASS CORE ;
    FOREIGN OA31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.430 3.285 0.620 ;
        RECT  3.155 1.040 3.265 1.470 ;
        RECT  3.050 1.040 3.155 1.150 ;
        RECT  2.750 0.430 3.050 1.150 ;
        RECT  2.625 0.430 2.750 0.620 ;
        RECT  2.745 1.040 2.750 1.150 ;
        RECT  2.635 1.040 2.745 1.470 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.900 2.150 1.100 ;
        RECT  1.850 0.760 1.950 1.100 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.900 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.710 1.350 0.900 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  0.550 1.010 1.050 1.100 ;
        RECT  0.450 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.710 1.625 0.960 ;
        RECT  1.450 0.710 1.550 1.300 ;
        RECT  0.360 1.210 1.450 1.300 ;
        RECT  0.270 1.020 0.360 1.300 ;
        RECT  0.170 1.020 0.270 1.120 ;
        RECT  0.050 0.680 0.170 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 -0.165 3.600 0.165 ;
        RECT  3.415 -0.165 3.525 0.695 ;
        RECT  0.000 -0.165 3.415 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 1.635 3.600 1.965 ;
        RECT  3.415 1.040 3.525 1.965 ;
        RECT  3.015 1.635 3.415 1.965 ;
        RECT  2.885 1.260 3.015 1.965 ;
        RECT  2.370 1.635 2.885 1.965 ;
        RECT  2.370 1.390 2.535 1.490 ;
        RECT  2.230 1.390 2.370 1.965 ;
        RECT  2.120 1.390 2.230 1.490 ;
        RECT  0.180 1.635 2.230 1.965 ;
        RECT  0.060 1.230 0.180 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 0.430 3.285 0.620 ;
        RECT  3.155 1.040 3.265 1.470 ;
        RECT  3.150 1.040 3.155 1.150 ;
        RECT  2.625 0.430 2.650 0.620 ;
        RECT  2.635 1.040 2.650 1.470 ;
        RECT  2.415 0.780 2.640 0.890 ;
        RECT  2.315 0.500 2.415 1.300 ;
        RECT  0.200 0.310 2.325 0.410 ;
        RECT  0.310 0.500 2.315 0.600 ;
        RECT  1.815 1.210 2.315 1.300 ;
        RECT  1.725 1.210 1.815 1.490 ;
        RECT  0.810 1.390 1.725 1.490 ;
        RECT  0.090 0.310 0.200 0.560 ;
    END
END OA31D4

MACRO OA32D0
    CLASS CORE ;
    FOREIGN OA32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.320 1.950 1.490 ;
        RECT  1.750 0.320 1.850 0.440 ;
        RECT  1.810 1.320 1.850 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.685 0.550 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.890 0.770 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.150 1.290 ;
        RECT  0.990 0.910 1.040 1.080 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.890 1.360 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.640 -0.165 2.000 0.165 ;
        RECT  1.500 -0.165 1.640 0.480 ;
        RECT  0.000 -0.165 1.500 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 1.635 2.000 1.965 ;
        RECT  0.065 1.295 0.195 1.965 ;
        RECT  0.000 1.635 0.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.580 0.650 1.700 1.490 ;
        RECT  0.825 0.650 1.580 0.775 ;
        RECT  0.560 1.385 1.580 1.490 ;
        RECT  0.085 0.300 1.280 0.470 ;
    END
END OA32D0

MACRO OA32D1
    CLASS CORE ;
    FOREIGN OA32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.295 2.150 1.490 ;
        RECT  2.005 0.295 2.050 0.675 ;
        RECT  2.005 1.265 2.050 1.490 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.160 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.090 ;
        RECT  1.340 0.700 1.450 0.910 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.820 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.855 -0.165 2.200 0.165 ;
        RECT  1.745 -0.165 1.855 0.665 ;
        RECT  0.000 -0.165 1.745 0.165 ;
        RECT  1.075 0.500 1.745 0.590 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.635 2.200 1.965 ;
        RECT  1.770 1.390 1.895 1.495 ;
        RECT  1.630 1.390 1.770 1.965 ;
        RECT  1.365 1.390 1.630 1.495 ;
        RECT  0.235 1.635 1.630 1.965 ;
        RECT  0.055 1.390 0.235 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.830 0.775 1.940 1.120 ;
        RECT  1.815 1.030 1.830 1.120 ;
        RECT  1.715 1.030 1.815 1.300 ;
        RECT  0.350 1.210 1.715 1.300 ;
        RECT  0.295 0.310 1.580 0.410 ;
        RECT  0.350 0.500 0.755 0.590 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.075 0.350 0.185 0.590 ;
    END
END OA32D1

MACRO OA32D2
    CLASS CORE ;
    FOREIGN OA32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.585 2.150 1.150 ;
        RECT  2.050 0.275 2.065 1.470 ;
        RECT  1.955 0.275 2.050 0.695 ;
        RECT  1.955 1.040 2.050 1.470 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.160 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.090 ;
        RECT  1.340 0.700 1.450 0.910 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.820 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 -0.165 2.400 0.165 ;
        RECT  2.215 -0.165 2.325 0.475 ;
        RECT  1.805 -0.165 2.215 0.165 ;
        RECT  1.695 -0.165 1.805 0.695 ;
        RECT  0.000 -0.165 1.695 0.165 ;
        RECT  1.075 0.500 1.695 0.590 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 1.635 2.400 1.965 ;
        RECT  2.215 1.260 2.325 1.965 ;
        RECT  1.770 1.635 2.215 1.965 ;
        RECT  1.770 1.390 1.845 1.495 ;
        RECT  1.635 1.390 1.770 1.965 ;
        RECT  1.365 1.390 1.635 1.495 ;
        RECT  0.235 1.635 1.635 1.965 ;
        RECT  0.055 1.390 0.235 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.815 0.805 1.940 0.915 ;
        RECT  1.715 0.805 1.815 1.300 ;
        RECT  0.350 1.210 1.715 1.300 ;
        RECT  0.295 0.310 1.575 0.410 ;
        RECT  0.350 0.500 0.755 0.590 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.075 0.350 0.185 0.590 ;
    END
END OA32D2

MACRO OA32D4
    CLASS CORE ;
    FOREIGN OA32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.755 0.275 3.865 0.695 ;
        RECT  3.755 1.040 3.865 1.470 ;
        RECT  3.650 0.585 3.755 0.695 ;
        RECT  3.650 1.040 3.755 1.150 ;
        RECT  3.350 0.585 3.650 1.150 ;
        RECT  3.345 0.585 3.350 0.695 ;
        RECT  3.345 1.040 3.350 1.150 ;
        RECT  3.235 0.275 3.345 0.695 ;
        RECT  3.235 1.040 3.345 1.470 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.420 0.910 2.550 1.090 ;
        RECT  2.250 0.790 2.420 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.645 0.590 2.750 1.090 ;
        RECT  1.985 0.590 2.645 0.680 ;
        RECT  1.885 0.590 1.985 0.960 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.710 1.350 1.090 ;
        RECT  0.550 1.000 1.225 1.090 ;
        RECT  0.450 0.710 0.550 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.775 1.605 0.965 ;
        RECT  1.450 0.775 1.550 1.290 ;
        RECT  0.360 1.200 1.450 1.290 ;
        RECT  0.270 1.020 0.360 1.290 ;
        RECT  0.170 1.020 0.270 1.120 ;
        RECT  0.050 0.710 0.170 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.695 ;
        RECT  3.605 -0.165 4.015 0.165 ;
        RECT  3.495 -0.165 3.605 0.475 ;
        RECT  2.100 -0.165 3.495 0.165 ;
        RECT  1.910 -0.165 2.100 0.300 ;
        RECT  0.000 -0.165 1.910 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.040 4.125 1.965 ;
        RECT  3.605 1.635 4.015 1.965 ;
        RECT  3.495 1.260 3.605 1.965 ;
        RECT  2.960 1.635 3.495 1.965 ;
        RECT  2.960 1.390 3.125 1.490 ;
        RECT  2.850 1.390 2.960 1.965 ;
        RECT  2.680 1.390 2.850 1.490 ;
        RECT  0.180 1.635 2.850 1.965 ;
        RECT  0.075 1.230 0.180 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.755 0.275 3.865 0.695 ;
        RECT  3.755 1.040 3.865 1.470 ;
        RECT  3.750 0.585 3.755 0.695 ;
        RECT  3.750 1.040 3.755 1.150 ;
        RECT  3.235 0.275 3.250 0.695 ;
        RECT  3.235 1.040 3.250 1.470 ;
        RECT  3.000 0.785 3.240 0.890 ;
        RECT  2.900 0.785 3.000 1.300 ;
        RECT  1.795 1.210 2.900 1.300 ;
        RECT  1.805 0.390 2.890 0.480 ;
        RECT  1.650 0.310 1.805 0.480 ;
        RECT  1.695 0.570 1.795 1.490 ;
        RECT  1.540 0.570 1.695 0.660 ;
        RECT  0.810 1.380 1.695 1.490 ;
        RECT  0.200 0.310 1.650 0.410 ;
        RECT  1.450 0.500 1.540 0.660 ;
        RECT  0.310 0.500 1.450 0.600 ;
        RECT  0.090 0.310 0.200 0.560 ;
    END
END OA32D4

MACRO OA33D0
    CLASS CORE ;
    FOREIGN OA33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.295 2.150 1.505 ;
        RECT  2.005 0.295 2.050 0.485 ;
        RECT  1.975 1.415 2.050 1.505 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  1.000 0.710 1.050 0.930 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.710 1.450 0.930 ;
        RECT  1.250 0.710 1.350 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.560 0.710 1.650 0.930 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.930 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.555 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.850 -0.165 2.200 0.165 ;
        RECT  1.740 -0.165 1.850 0.600 ;
        RECT  0.000 -0.165 1.740 0.165 ;
        RECT  1.140 0.500 1.740 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.865 1.635 2.200 1.965 ;
        RECT  1.670 1.415 1.865 1.965 ;
        RECT  0.235 1.635 1.670 1.965 ;
        RECT  0.055 1.410 0.235 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.870 0.775 1.960 1.305 ;
        RECT  1.030 1.200 1.870 1.305 ;
        RECT  0.285 0.300 1.635 0.410 ;
        RECT  0.850 1.200 1.030 1.510 ;
        RECT  0.350 1.200 0.850 1.310 ;
        RECT  0.350 0.500 0.780 0.600 ;
        RECT  0.260 0.500 0.350 1.310 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.075 0.280 0.185 0.590 ;
    END
END OA33D0

MACRO OA33D1
    CLASS CORE ;
    FOREIGN OA33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.295 2.150 1.505 ;
        RECT  2.005 0.295 2.050 0.675 ;
        RECT  1.975 1.415 2.050 1.505 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.980 0.710 1.050 0.930 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.710 1.450 0.930 ;
        RECT  1.250 0.710 1.350 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.560 0.710 1.650 0.930 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.930 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.555 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.825 -0.165 2.200 0.165 ;
        RECT  1.715 -0.165 1.825 0.600 ;
        RECT  0.000 -0.165 1.715 0.165 ;
        RECT  1.075 0.500 1.715 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.865 1.635 2.200 1.965 ;
        RECT  1.660 1.400 1.865 1.965 ;
        RECT  0.235 1.635 1.660 1.965 ;
        RECT  0.055 1.410 0.235 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.870 0.775 1.960 1.290 ;
        RECT  0.350 1.200 1.870 1.290 ;
        RECT  0.295 0.310 1.580 0.410 ;
        RECT  0.350 0.500 0.755 0.600 ;
        RECT  0.260 0.500 0.350 1.290 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.060 0.350 0.185 0.590 ;
    END
END OA33D1

MACRO OA33D2
    CLASS CORE ;
    FOREIGN OA33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.555 2.150 1.160 ;
        RECT  2.050 0.555 2.130 1.500 ;
        RECT  1.940 0.295 2.050 0.665 ;
        RECT  2.040 1.040 2.050 1.500 ;
        RECT  1.910 1.390 2.040 1.500 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.980 0.710 1.050 0.930 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.710 1.430 0.930 ;
        RECT  1.250 0.710 1.350 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.585 0.710 1.650 0.930 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.930 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.555 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 -0.165 2.400 0.165 ;
        RECT  2.205 -0.165 2.315 0.445 ;
        RECT  1.790 -0.165 2.205 0.165 ;
        RECT  1.680 -0.165 1.790 0.600 ;
        RECT  0.000 -0.165 1.680 0.165 ;
        RECT  1.075 0.500 1.680 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.635 2.400 1.965 ;
        RECT  2.225 1.355 2.320 1.965 ;
        RECT  1.820 1.635 2.225 1.965 ;
        RECT  1.645 1.390 1.820 1.965 ;
        RECT  0.235 1.635 1.645 1.965 ;
        RECT  0.055 1.390 0.235 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.860 0.775 1.950 1.300 ;
        RECT  0.350 1.200 1.860 1.300 ;
        RECT  0.295 0.310 1.570 0.410 ;
        RECT  0.350 0.500 0.745 0.600 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.060 0.350 0.185 0.590 ;
    END
END OA33D2

MACRO OA33D4
    CLASS CORE ;
    FOREIGN OA33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.155 0.275 4.265 0.695 ;
        RECT  4.155 1.045 4.265 1.475 ;
        RECT  4.050 0.585 4.155 0.695 ;
        RECT  4.050 1.045 4.155 1.155 ;
        RECT  3.750 0.585 4.050 1.155 ;
        RECT  3.745 0.585 3.750 0.695 ;
        RECT  3.745 1.045 3.750 1.155 ;
        RECT  3.635 0.275 3.745 0.695 ;
        RECT  3.635 1.045 3.745 1.475 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1104 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.710 1.350 0.900 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.550 1.000 1.050 1.090 ;
        RECT  0.450 0.700 0.550 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1101 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.710 1.560 1.290 ;
        RECT  0.360 1.200 1.440 1.290 ;
        RECT  0.270 1.020 0.360 1.290 ;
        RECT  0.170 1.020 0.270 1.120 ;
        RECT  0.050 0.680 0.170 1.120 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.550 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.805 0.710 2.950 1.090 ;
        RECT  2.150 1.000 2.805 1.090 ;
        RECT  1.985 0.710 2.150 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1093 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.045 0.710 3.160 1.290 ;
        RECT  1.805 1.200 3.045 1.290 ;
        RECT  1.650 0.710 1.805 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 -0.165 4.600 0.165 ;
        RECT  4.415 -0.165 4.525 0.695 ;
        RECT  4.005 -0.165 4.415 0.165 ;
        RECT  3.895 -0.165 4.005 0.475 ;
        RECT  0.000 -0.165 3.895 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.635 4.600 1.965 ;
        RECT  4.415 1.045 4.525 1.965 ;
        RECT  4.005 1.635 4.415 1.965 ;
        RECT  3.895 1.265 4.005 1.965 ;
        RECT  0.180 1.635 3.895 1.965 ;
        RECT  0.060 1.230 0.180 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.155 0.275 4.265 0.695 ;
        RECT  4.155 1.045 4.265 1.475 ;
        RECT  4.150 0.585 4.155 0.695 ;
        RECT  4.150 1.045 4.155 1.155 ;
        RECT  3.635 0.275 3.650 0.695 ;
        RECT  3.635 1.045 3.650 1.475 ;
        RECT  3.370 0.785 3.595 0.900 ;
        RECT  3.270 0.500 3.370 1.500 ;
        RECT  0.195 0.310 3.300 0.410 ;
        RECT  1.800 0.500 3.270 0.600 ;
        RECT  0.800 1.400 3.270 1.500 ;
        RECT  0.075 0.310 0.195 0.560 ;
    END
END OA33D4

MACRO OAI211D0
    CLASS CORE ;
    FOREIGN OAI211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1420 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.300 ;
        RECT  0.310 0.500 1.250 0.600 ;
        RECT  0.945 1.210 1.250 1.300 ;
        RECT  0.835 1.210 0.945 1.490 ;
        RECT  0.185 1.210 0.835 1.300 ;
        RECT  0.075 1.210 0.185 1.490 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.930 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.850 0.930 ;
        RECT  0.650 0.710 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.560 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.165 1.400 0.165 ;
        RECT  1.150 -0.165 1.320 0.390 ;
        RECT  0.000 -0.165 1.150 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.635 1.400 1.965 ;
        RECT  1.090 1.410 1.260 1.965 ;
        RECT  0.690 1.635 1.090 1.965 ;
        RECT  0.520 1.410 0.690 1.965 ;
        RECT  0.000 1.635 0.520 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.185 0.300 0.805 0.410 ;
        RECT  0.075 0.300 0.185 0.500 ;
    END
END OAI211D0

MACRO OAI211D1
    CLASS CORE ;
    FOREIGN OAI211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2650 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.300 ;
        RECT  0.305 0.500 1.250 0.590 ;
        RECT  0.045 1.210 1.250 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.970 0.700 1.050 0.950 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.165 1.400 0.165 ;
        RECT  1.050 -0.165 1.220 0.390 ;
        RECT  0.000 -0.165 1.050 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.635 1.400 1.965 ;
        RECT  1.090 1.410 1.260 1.965 ;
        RECT  0.690 1.635 1.090 1.965 ;
        RECT  0.520 1.410 0.690 1.965 ;
        RECT  0.000 1.635 0.520 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.190 0.310 0.755 0.410 ;
        RECT  0.070 0.310 0.190 0.560 ;
    END
END OAI211D1

MACRO OAI211D2
    CLASS CORE ;
    FOREIGN OAI211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 2.350 1.295 ;
        RECT  1.340 0.510 2.250 0.600 ;
        RECT  0.300 1.200 2.250 1.295 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.710 1.150 1.090 ;
        RECT  0.170 1.000 1.030 1.090 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.950 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1093 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.710 2.150 1.090 ;
        RECT  1.370 1.000 2.050 1.090 ;
        RECT  1.250 0.710 1.370 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.165 2.400 0.165 ;
        RECT  0.565 -0.165 0.745 0.410 ;
        RECT  0.000 -0.165 0.565 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.335 1.635 2.400 1.965 ;
        RECT  2.165 1.405 2.335 1.965 ;
        RECT  0.970 1.635 2.165 1.965 ;
        RECT  0.970 1.390 1.280 1.490 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.550 1.390 0.830 1.490 ;
        RECT  0.190 1.635 0.830 1.965 ;
        RECT  0.080 1.240 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.230 0.300 2.335 0.400 ;
        RECT  1.120 0.300 1.230 0.590 ;
        RECT  0.190 0.500 1.120 0.590 ;
        RECT  0.065 0.350 0.190 0.590 ;
    END
END OAI211D2

MACRO OAI211D4
    CLASS CORE ;
    FOREIGN OAI211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9980 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.210 4.460 1.300 ;
        RECT  2.650 0.950 2.750 1.300 ;
        RECT  2.350 0.950 2.650 1.050 ;
        RECT  2.250 0.500 2.350 1.050 ;
        RECT  1.050 0.500 2.250 0.590 ;
        RECT  0.750 0.500 1.050 1.300 ;
        RECT  0.070 0.500 0.750 0.590 ;
        RECT  0.340 1.210 0.750 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.700 4.155 1.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.045 0.700 3.155 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.700 0.555 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.700 1.955 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 -0.165 4.800 0.165 ;
        RECT  4.170 0.310 4.470 0.410 ;
        RECT  4.030 -0.165 4.170 0.410 ;
        RECT  0.000 -0.165 4.030 0.165 ;
        RECT  3.740 0.310 4.030 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 1.635 4.800 1.965 ;
        RECT  4.170 1.390 4.730 1.490 ;
        RECT  4.030 1.390 4.170 1.965 ;
        RECT  3.480 1.390 4.030 1.490 ;
        RECT  2.970 1.635 4.030 1.965 ;
        RECT  2.970 1.390 3.170 1.490 ;
        RECT  2.830 1.390 2.970 1.965 ;
        RECT  2.440 1.390 2.830 1.490 ;
        RECT  1.770 1.635 2.830 1.965 ;
        RECT  1.770 1.390 2.130 1.490 ;
        RECT  1.630 1.390 1.770 1.965 ;
        RECT  1.400 1.390 1.630 1.490 ;
        RECT  0.000 1.635 1.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 1.210 4.460 1.300 ;
        RECT  2.650 0.950 2.750 1.300 ;
        RECT  2.350 0.950 2.650 1.050 ;
        RECT  2.250 0.500 2.350 1.050 ;
        RECT  1.150 0.500 2.250 0.590 ;
        RECT  0.070 0.500 0.650 0.590 ;
        RECT  0.340 1.210 0.650 1.300 ;
        RECT  2.460 0.500 4.730 0.590 ;
        RECT  0.340 0.310 3.420 0.410 ;
        RECT  1.270 1.210 2.380 1.300 ;
        RECT  1.160 1.210 1.270 1.490 ;
        RECT  0.225 1.390 1.160 1.490 ;
        RECT  0.105 1.030 0.225 1.490 ;
    END
END OAI211D4

MACRO OAI21D0
    CLASS CORE ;
    FOREIGN OAI21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.500 1.150 1.340 ;
        RECT  0.310 0.500 1.035 0.600 ;
        RECT  0.715 1.240 1.035 1.340 ;
        RECT  0.605 1.240 0.715 1.490 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.850 0.970 ;
        RECT  0.650 0.710 0.750 1.120 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.165 1.200 0.165 ;
        RECT  0.915 -0.165 1.070 0.390 ;
        RECT  0.000 -0.165 0.915 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.635 1.200 1.965 ;
        RECT  0.860 1.455 1.030 1.965 ;
        RECT  0.190 1.635 0.860 1.965 ;
        RECT  0.070 1.325 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.185 0.300 0.805 0.410 ;
        RECT  0.075 0.300 0.185 0.500 ;
    END
END OAI21D0

MACRO OAI21D1
    CLASS CORE ;
    FOREIGN OAI21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.500 1.150 1.340 ;
        RECT  0.305 0.500 1.050 0.590 ;
        RECT  0.555 1.240 1.050 1.340 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.970 ;
        RECT  0.650 0.700 0.750 1.120 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.550 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.165 1.200 0.165 ;
        RECT  0.875 -0.165 1.030 0.390 ;
        RECT  0.000 -0.165 0.875 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.635 1.200 1.965 ;
        RECT  0.860 1.450 1.030 1.965 ;
        RECT  0.190 1.635 0.860 1.965 ;
        RECT  0.070 1.325 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.195 0.310 0.765 0.410 ;
        RECT  0.070 0.310 0.195 0.560 ;
    END
END OAI21D1

MACRO OAI21D2
    CLASS CORE ;
    FOREIGN OAI21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4260 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.210 1.750 1.490 ;
        RECT  0.550 1.210 1.615 1.300 ;
        RECT  0.550 0.500 1.505 0.590 ;
        RECT  0.450 0.500 0.550 1.300 ;
        RECT  0.185 1.210 0.450 1.300 ;
        RECT  0.050 1.210 0.185 1.490 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.700 0.360 1.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.700 1.150 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.700 1.550 1.100 ;
        RECT  0.760 1.010 1.440 1.100 ;
        RECT  0.645 0.700 0.760 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.245 1.635 1.800 1.965 ;
        RECT  1.065 1.390 1.245 1.965 ;
        RECT  0.000 1.635 1.065 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.615 0.310 1.725 0.585 ;
        RECT  0.185 0.310 1.615 0.410 ;
        RECT  0.075 0.310 0.185 0.570 ;
    END
END OAI21D2

MACRO OAI21D4
    CLASS CORE ;
    FOREIGN OAI21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 1.210 3.305 1.300 ;
        RECT  2.535 0.500 2.635 1.300 ;
        RECT  0.650 0.500 2.535 0.600 ;
        RECT  0.650 1.200 1.005 1.300 ;
        RECT  0.350 0.500 0.650 1.300 ;
        RECT  0.045 0.500 0.350 0.600 ;
        RECT  0.295 1.200 0.350 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.795 0.710 3.205 0.890 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.395 0.710 2.205 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 0.710 1.155 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.635 3.600 1.965 ;
        RECT  2.970 1.390 3.555 1.500 ;
        RECT  2.830 1.390 2.970 1.965 ;
        RECT  2.325 1.390 2.830 1.500 ;
        RECT  1.770 1.635 2.830 1.965 ;
        RECT  1.770 1.390 2.015 1.500 ;
        RECT  1.630 1.390 1.770 1.965 ;
        RECT  1.305 1.390 1.630 1.500 ;
        RECT  0.000 1.635 1.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.635 1.210 3.305 1.300 ;
        RECT  2.535 0.500 2.635 1.300 ;
        RECT  0.750 0.500 2.535 0.600 ;
        RECT  0.750 1.200 1.005 1.300 ;
        RECT  0.045 0.500 0.250 0.600 ;
        RECT  0.285 0.300 3.555 0.410 ;
        RECT  1.655 1.210 2.265 1.300 ;
        RECT  1.545 1.000 1.655 1.300 ;
        RECT  1.215 1.000 1.545 1.090 ;
        RECT  1.115 1.000 1.215 1.490 ;
        RECT  0.185 1.390 1.115 1.490 ;
        RECT  0.075 1.020 0.185 1.490 ;
    END
END OAI21D4

MACRO OAI221D0
    CLASS CORE ;
    FOREIGN OAI221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1430 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.410 1.530 1.520 ;
        RECT  0.865 0.495 0.995 0.730 ;
        RECT  0.150 0.495 0.865 0.585 ;
        RECT  0.050 0.495 0.150 1.520 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.350 1.290 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.555 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.595 1.550 1.300 ;
        RECT  0.840 1.210 1.440 1.300 ;
        RECT  0.650 1.070 0.840 1.300 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.870 1.150 1.105 ;
        RECT  0.775 0.870 0.960 0.960 ;
        RECT  0.650 0.695 0.775 0.960 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.680 1.350 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.600 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.405 0.275 1.535 0.480 ;
        RECT  0.285 0.275 1.405 0.405 ;
    END
END OAI221D0

MACRO OAI221D1
    CLASS CORE ;
    FOREIGN OAI221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.200 1.515 1.290 ;
        RECT  0.150 0.510 0.495 0.600 ;
        RECT  0.050 0.510 0.150 1.290 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.580 0.710 1.650 0.930 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 0.710 1.380 0.930 ;
        RECT  1.250 0.710 1.360 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.940 0.805 1.150 1.090 ;
        RECT  0.850 0.910 0.940 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.355 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.710 0.610 0.930 ;
        RECT  0.450 0.710 0.560 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.585 ;
        RECT  0.000 -0.165 1.615 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.635 1.800 1.965 ;
        RECT  1.615 1.200 1.725 1.965 ;
        RECT  0.760 1.635 1.615 1.965 ;
        RECT  0.760 1.390 1.015 1.500 ;
        RECT  0.630 1.390 0.760 1.965 ;
        RECT  0.045 1.400 0.630 1.510 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.945 0.500 1.515 0.600 ;
        RECT  0.045 0.290 1.255 0.400 ;
        RECT  0.835 0.500 0.945 0.705 ;
    END
END OAI221D1

MACRO OAI221D2
    CLASS CORE ;
    FOREIGN OAI221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.500 3.150 1.300 ;
        RECT  1.900 0.500 3.050 0.600 ;
        RECT  0.050 1.200 3.050 1.300 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.360 1.090 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  0.950 1.000 1.650 1.090 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.765 0.710 0.850 0.920 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.750 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 2.950 1.090 ;
        RECT  2.150 1.000 2.850 1.090 ;
        RECT  2.040 0.710 2.150 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.165 3.200 0.165 ;
        RECT  0.305 -0.165 0.485 0.410 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.605 1.635 3.200 1.965 ;
        RECT  2.425 1.390 2.605 1.965 ;
        RECT  0.770 1.635 2.425 1.965 ;
        RECT  0.770 1.390 1.280 1.500 ;
        RECT  0.630 1.390 0.770 1.965 ;
        RECT  0.290 1.390 0.630 1.500 ;
        RECT  0.000 1.635 0.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.810 0.300 2.880 0.410 ;
        RECT  0.185 0.500 1.790 0.600 ;
        RECT  0.065 0.350 0.185 0.600 ;
    END
END OAI221D2

MACRO OAI221D4
    CLASS CORE ;
    FOREIGN OAI221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.275 3.065 0.695 ;
        RECT  2.955 1.040 3.065 1.470 ;
        RECT  2.850 0.585 2.955 0.695 ;
        RECT  2.850 1.040 2.955 1.150 ;
        RECT  2.550 0.585 2.850 1.150 ;
        RECT  2.545 0.585 2.550 0.695 ;
        RECT  2.545 1.040 2.550 1.150 ;
        RECT  2.435 0.275 2.545 0.695 ;
        RECT  2.435 1.040 2.545 1.470 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.700 1.600 0.950 ;
        RECT  1.450 0.700 1.550 1.100 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.355 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.700 0.950 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.570 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 -0.165 3.400 0.165 ;
        RECT  3.210 -0.165 3.330 0.695 ;
        RECT  2.805 -0.165 3.210 0.165 ;
        RECT  2.695 -0.165 2.805 0.475 ;
        RECT  2.290 -0.165 2.695 0.165 ;
        RECT  2.170 -0.165 2.290 0.695 ;
        RECT  1.765 -0.165 2.170 0.165 ;
        RECT  1.655 -0.165 1.765 0.585 ;
        RECT  0.000 -0.165 1.655 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 1.635 3.400 1.965 ;
        RECT  3.210 1.040 3.330 1.965 ;
        RECT  2.805 1.635 3.210 1.965 ;
        RECT  2.695 1.260 2.805 1.965 ;
        RECT  2.290 1.635 2.695 1.965 ;
        RECT  2.170 1.040 2.290 1.965 ;
        RECT  0.970 1.635 2.170 1.965 ;
        RECT  0.970 1.390 1.805 1.500 ;
        RECT  0.835 1.390 0.970 1.965 ;
        RECT  0.055 1.390 0.835 1.500 ;
        RECT  0.000 1.635 0.835 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.955 0.275 3.065 0.695 ;
        RECT  2.955 1.040 3.065 1.470 ;
        RECT  2.950 0.585 2.955 0.695 ;
        RECT  2.950 1.040 2.955 1.150 ;
        RECT  2.435 0.275 2.450 0.695 ;
        RECT  2.435 1.040 2.450 1.470 ;
        RECT  2.060 0.785 2.430 0.890 ;
        RECT  1.960 0.275 2.060 1.475 ;
        RECT  1.920 0.275 1.960 0.675 ;
        RECT  1.920 1.045 1.960 1.475 ;
        RECT  1.810 0.775 1.850 0.945 ;
        RECT  1.710 0.775 1.810 1.300 ;
        RECT  0.360 1.210 1.710 1.300 ;
        RECT  0.825 0.500 1.545 0.590 ;
        RECT  0.715 0.300 1.295 0.410 ;
        RECT  0.605 0.300 0.715 0.590 ;
        RECT  0.180 0.300 0.605 0.390 ;
        RECT  0.360 0.500 0.505 0.590 ;
        RECT  0.270 0.500 0.360 1.300 ;
        RECT  0.060 0.300 0.180 0.560 ;
    END
END OAI221D4

MACRO OAI221XD4
    CLASS CORE ;
    FOREIGN OAI221XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.500 5.695 0.600 ;
        RECT  4.250 1.000 4.655 1.115 ;
        RECT  3.950 0.500 4.250 1.115 ;
        RECT  3.935 0.500 3.950 0.600 ;
        RECT  0.965 1.000 3.950 1.115 ;
        RECT  0.855 1.000 0.965 1.470 ;
        RECT  0.445 1.000 0.855 1.110 ;
        RECT  0.335 1.000 0.445 1.470 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 3.150 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.710 5.550 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.710 4.750 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 -0.165 6.000 0.165 ;
        RECT  0.970 0.300 1.255 0.410 ;
        RECT  0.830 -0.165 0.970 0.410 ;
        RECT  0.185 -0.165 0.830 0.165 ;
        RECT  0.555 0.300 0.830 0.410 ;
        RECT  0.075 -0.165 0.185 0.695 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.645 1.635 6.000 1.965 ;
        RECT  5.535 1.260 5.645 1.965 ;
        RECT  5.125 1.635 5.535 1.965 ;
        RECT  5.015 1.260 5.125 1.965 ;
        RECT  1.970 1.635 5.015 1.965 ;
        RECT  1.970 1.395 2.315 1.505 ;
        RECT  1.830 1.395 1.970 1.965 ;
        RECT  1.585 1.395 1.830 1.505 ;
        RECT  1.225 1.635 1.830 1.965 ;
        RECT  1.115 1.235 1.225 1.965 ;
        RECT  0.705 1.635 1.115 1.965 ;
        RECT  0.595 1.235 0.705 1.965 ;
        RECT  0.185 1.635 0.595 1.965 ;
        RECT  0.075 1.040 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.350 0.500 5.695 0.600 ;
        RECT  4.350 1.000 4.655 1.115 ;
        RECT  0.965 1.000 3.850 1.115 ;
        RECT  0.855 1.000 0.965 1.470 ;
        RECT  0.445 1.000 0.855 1.110 ;
        RECT  0.335 1.000 0.445 1.470 ;
        RECT  3.825 0.300 5.945 0.410 ;
        RECT  5.795 1.040 5.905 1.470 ;
        RECT  5.385 1.040 5.795 1.150 ;
        RECT  5.275 1.040 5.385 1.470 ;
        RECT  4.865 1.040 5.275 1.150 ;
        RECT  4.755 1.040 4.865 1.470 ;
        RECT  3.685 1.370 4.755 1.470 ;
        RECT  3.715 0.300 3.825 0.695 ;
        RECT  3.565 0.300 3.715 0.410 ;
        RECT  1.335 1.205 3.595 1.305 ;
        RECT  3.455 0.300 3.565 0.695 ;
        RECT  1.345 0.300 3.455 0.410 ;
        RECT  0.445 0.520 3.345 0.620 ;
        RECT  0.335 0.275 0.445 0.695 ;
    END
END OAI221XD4

MACRO OAI222D0
    CLASS CORE ;
    FOREIGN OAI222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1430 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.410 1.730 1.520 ;
        RECT  1.070 0.495 1.195 0.730 ;
        RECT  0.430 0.495 1.070 0.585 ;
        RECT  0.340 0.495 0.430 0.655 ;
        RECT  0.150 0.565 0.340 0.655 ;
        RECT  0.050 0.565 0.150 1.520 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.765 0.560 1.290 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.765 0.350 1.290 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.755 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.595 1.750 1.300 ;
        RECT  1.040 1.210 1.640 1.300 ;
        RECT  0.850 1.070 1.040 1.300 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.870 1.350 1.105 ;
        RECT  0.980 0.870 1.160 0.960 ;
        RECT  0.850 0.695 0.980 0.960 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.680 1.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.605 0.275 1.735 0.480 ;
        RECT  0.200 0.275 1.605 0.405 ;
        RECT  0.060 0.275 0.200 0.445 ;
    END
END OAI222D0

MACRO OAI222D1
    CLASS CORE ;
    FOREIGN OAI222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2730 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.210 1.575 1.300 ;
        RECT  0.150 0.500 0.515 0.590 ;
        RECT  0.050 0.500 0.150 1.300 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.700 1.950 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.790 0.700 0.850 0.950 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.160 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.360 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.605 0.950 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 -0.165 2.200 0.165 ;
        RECT  1.945 -0.165 2.055 0.585 ;
        RECT  1.510 -0.165 1.945 0.165 ;
        RECT  1.510 0.300 1.585 0.410 ;
        RECT  1.395 -0.165 1.510 0.410 ;
        RECT  0.000 -0.165 1.395 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.005 1.635 2.200 1.965 ;
        RECT  1.895 1.210 2.005 1.965 ;
        RECT  1.205 1.635 1.895 1.965 ;
        RECT  1.205 1.390 1.295 1.500 ;
        RECT  1.095 1.390 1.205 1.965 ;
        RECT  0.165 1.635 1.095 1.965 ;
        RECT  0.165 1.410 0.265 1.520 ;
        RECT  0.055 1.410 0.165 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.845 0.500 1.835 0.590 ;
        RECT  0.050 0.285 1.285 0.390 ;
    END
END OAI222D1

MACRO OAI222D2
    CLASS CORE ;
    FOREIGN OAI222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5810 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.295 3.555 1.300 ;
        RECT  2.345 0.295 3.450 0.405 ;
        RECT  0.525 1.200 3.450 1.300 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.710 1.150 1.090 ;
        RECT  0.170 1.000 0.995 1.090 ;
        RECT  0.050 0.710 0.170 1.090 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.710 2.150 1.090 ;
        RECT  1.350 1.000 2.040 1.090 ;
        RECT  1.240 0.710 1.350 1.090 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 3.150 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.710 3.360 1.090 ;
        RECT  2.555 1.000 3.250 1.090 ;
        RECT  2.445 0.710 2.555 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.635 3.600 1.965 ;
        RECT  2.370 1.390 3.055 1.500 ;
        RECT  2.230 1.390 2.370 1.965 ;
        RECT  1.025 1.390 2.230 1.500 ;
        RECT  0.190 1.635 2.230 1.965 ;
        RECT  0.070 1.240 0.190 1.965 ;
        RECT  0.000 1.635 0.070 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.285 0.495 3.315 0.600 ;
        RECT  0.045 0.295 2.255 0.405 ;
    END
END OAI222D2

MACRO OAI222D4
    CLASS CORE ;
    FOREIGN OAI222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.545 2.840 0.720 ;
        RECT  2.450 1.230 2.840 1.470 ;
        RECT  2.130 0.545 2.450 1.470 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.700 1.555 1.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.700 1.830 0.910 ;
        RECT  1.650 0.700 1.750 1.100 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.805 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.700 1.155 1.100 ;
        RECT  0.975 0.700 1.045 0.910 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.050 1.635 3.400 1.965 ;
        RECT  2.940 1.255 3.050 1.965 ;
        RECT  2.040 1.635 2.940 1.965 ;
        RECT  1.870 1.395 2.040 1.965 ;
        RECT  1.240 1.635 1.870 1.965 ;
        RECT  1.070 1.390 1.240 1.965 ;
        RECT  0.280 1.635 1.070 1.965 ;
        RECT  0.090 1.390 0.280 1.965 ;
        RECT  0.000 1.635 0.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.545 2.840 0.720 ;
        RECT  2.550 1.230 2.840 1.470 ;
        RECT  3.250 0.285 3.350 1.490 ;
        RECT  3.210 0.285 3.250 0.675 ;
        RECT  3.210 1.030 3.250 1.490 ;
        RECT  2.920 1.030 3.210 1.120 ;
        RECT  3.100 0.765 3.130 0.935 ;
        RECT  3.010 0.360 3.100 0.935 ;
        RECT  2.020 0.360 3.010 0.450 ;
        RECT  2.830 0.810 2.920 1.120 ;
        RECT  2.610 0.810 2.830 0.920 ;
        RECT  1.930 0.360 2.020 1.300 ;
        RECT  0.360 1.210 1.930 1.300 ;
        RECT  0.820 0.500 1.800 0.590 ;
        RECT  0.060 0.300 1.270 0.410 ;
        RECT  0.360 0.500 0.510 0.590 ;
        RECT  0.260 0.500 0.360 1.300 ;
    END
END OAI222D4

MACRO OAI222XD4
    CLASS CORE ;
    FOREIGN OAI222XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.500 6.715 0.600 ;
        RECT  5.250 1.000 5.675 1.115 ;
        RECT  4.950 0.500 5.250 1.115 ;
        RECT  1.305 1.000 4.950 1.115 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.950 0.890 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.2197 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 3.150 0.890 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.710 6.550 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.710 5.750 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.970 -0.165 7.000 0.165 ;
        RECT  1.970 0.300 2.275 0.410 ;
        RECT  1.830 -0.165 1.970 0.410 ;
        RECT  1.255 -0.165 1.830 0.165 ;
        RECT  1.565 0.300 1.830 0.410 ;
        RECT  1.145 -0.165 1.255 0.410 ;
        RECT  0.185 -0.165 1.145 0.165 ;
        RECT  1.045 0.300 1.145 0.410 ;
        RECT  0.075 -0.165 0.185 0.695 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 1.635 7.000 1.965 ;
        RECT  6.555 1.260 6.665 1.965 ;
        RECT  6.145 1.635 6.555 1.965 ;
        RECT  6.035 1.260 6.145 1.965 ;
        RECT  2.970 1.635 6.035 1.965 ;
        RECT  2.970 1.395 3.335 1.505 ;
        RECT  2.830 1.395 2.970 1.965 ;
        RECT  2.605 1.395 2.830 1.505 ;
        RECT  0.445 1.635 2.830 1.965 ;
        RECT  0.335 1.260 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.350 0.500 6.715 0.600 ;
        RECT  5.350 1.000 5.675 1.115 ;
        RECT  1.305 1.000 4.850 1.115 ;
        RECT  6.825 0.300 6.935 0.510 ;
        RECT  6.815 1.040 6.925 1.470 ;
        RECT  4.840 0.300 6.825 0.410 ;
        RECT  6.405 1.040 6.815 1.150 ;
        RECT  6.295 1.040 6.405 1.470 ;
        RECT  5.885 1.040 6.295 1.150 ;
        RECT  5.775 1.040 5.885 1.470 ;
        RECT  4.705 1.370 5.775 1.470 ;
        RECT  4.735 0.300 4.840 0.695 ;
        RECT  4.585 0.300 4.735 0.410 ;
        RECT  2.355 1.205 4.615 1.305 ;
        RECT  4.475 0.300 4.585 0.695 ;
        RECT  2.365 0.300 4.475 0.410 ;
        RECT  1.465 0.520 4.365 0.620 ;
        RECT  1.205 1.360 2.275 1.470 ;
        RECT  1.355 0.275 1.465 0.695 ;
        RECT  0.445 0.500 1.355 0.600 ;
        RECT  1.095 1.040 1.205 1.470 ;
        RECT  0.705 1.040 1.095 1.150 ;
        RECT  0.595 1.040 0.705 1.470 ;
        RECT  0.185 1.040 0.595 1.150 ;
        RECT  0.335 0.275 0.445 0.695 ;
        RECT  0.075 1.040 0.185 1.470 ;
    END
END OAI222XD4

MACRO OAI22D0
    CLASS CORE ;
    FOREIGN OAI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.350 1.345 ;
        RECT  0.855 0.510 1.250 0.600 ;
        RECT  0.050 1.235 1.250 1.345 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.550 1.120 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.120 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.940 ;
        RECT  0.650 0.710 0.750 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.150 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 -0.165 1.400 0.165 ;
        RECT  0.410 0.300 0.510 0.410 ;
        RECT  0.300 -0.165 0.410 0.410 ;
        RECT  0.000 -0.165 0.300 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.635 1.400 1.965 ;
        RECT  0.580 1.455 0.750 1.965 ;
        RECT  0.000 1.635 0.580 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.290 1.340 0.400 ;
        RECT  0.610 0.290 0.720 0.590 ;
        RECT  0.200 0.500 0.610 0.590 ;
        RECT  0.090 0.265 0.200 0.590 ;
    END
END OAI22D0

MACRO OAI22D1
    CLASS CORE ;
    FOREIGN OAI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2650 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.345 ;
        RECT  0.830 0.500 1.250 0.590 ;
        RECT  0.050 1.235 1.250 1.345 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.550 1.120 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.120 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.810 0.970 ;
        RECT  0.650 0.700 0.750 1.120 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.700 1.150 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 -0.165 1.400 0.165 ;
        RECT  0.310 -0.165 0.500 0.410 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.635 1.400 1.965 ;
        RECT  0.580 1.455 0.750 1.965 ;
        RECT  0.000 1.635 0.580 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.300 1.305 0.390 ;
        RECT  0.610 0.300 0.720 0.590 ;
        RECT  0.200 0.500 0.610 0.590 ;
        RECT  0.090 0.350 0.200 0.590 ;
    END
END OAI22D1

MACRO OAI22D2
    CLASS CORE ;
    FOREIGN OAI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.500 2.350 1.300 ;
        RECT  1.340 0.500 2.250 0.590 ;
        RECT  0.545 1.210 2.250 1.300 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.700 1.150 1.100 ;
        RECT  0.170 1.010 1.030 1.100 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.750 0.900 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.700 2.150 1.100 ;
        RECT  1.370 1.010 2.050 1.100 ;
        RECT  1.250 0.700 1.370 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.700 1.950 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.165 2.400 0.165 ;
        RECT  0.770 0.310 1.010 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.300 0.310 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.635 2.400 1.965 ;
        RECT  1.080 1.390 1.270 1.965 ;
        RECT  0.190 1.635 1.080 1.965 ;
        RECT  0.080 1.240 0.190 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 0.290 2.300 0.390 ;
        RECT  1.125 0.290 1.225 0.590 ;
        RECT  0.185 0.500 1.125 0.590 ;
        RECT  0.080 0.350 0.185 0.590 ;
    END
END OAI22D2

MACRO OAI22D4
    CLASS CORE ;
    FOREIGN OAI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.145 1.210 4.705 1.300 ;
        RECT  4.035 1.010 4.145 1.300 ;
        RECT  2.350 1.010 4.035 1.100 ;
        RECT  2.250 0.500 2.350 1.100 ;
        RECT  0.850 0.500 2.250 0.590 ;
        RECT  0.850 1.210 1.005 1.300 ;
        RECT  0.550 0.500 0.850 1.300 ;
        RECT  0.045 0.500 0.550 0.590 ;
        RECT  0.295 1.210 0.550 1.300 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.700 3.150 0.900 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.700 4.555 1.100 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.700 1.755 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.355 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 -0.165 5.000 0.165 ;
        RECT  4.820 -0.165 4.930 0.560 ;
        RECT  4.170 -0.165 4.820 0.165 ;
        RECT  4.170 0.310 4.455 0.410 ;
        RECT  4.030 -0.165 4.170 0.410 ;
        RECT  3.170 -0.165 4.030 0.165 ;
        RECT  3.725 0.310 4.030 0.410 ;
        RECT  3.170 0.310 3.385 0.410 ;
        RECT  3.030 -0.165 3.170 0.410 ;
        RECT  0.000 -0.165 3.030 0.165 ;
        RECT  2.665 0.310 3.030 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.635 5.000 1.965 ;
        RECT  3.370 1.390 3.635 1.490 ;
        RECT  3.230 1.390 3.370 1.965 ;
        RECT  2.915 1.390 3.230 1.490 ;
        RECT  2.555 1.635 3.230 1.965 ;
        RECT  2.445 1.210 2.555 1.965 ;
        RECT  1.770 1.635 2.445 1.965 ;
        RECT  1.770 1.390 2.085 1.490 ;
        RECT  1.630 1.390 1.770 1.965 ;
        RECT  1.365 1.390 1.630 1.490 ;
        RECT  0.000 1.635 1.630 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.145 1.210 4.705 1.300 ;
        RECT  4.035 1.010 4.145 1.300 ;
        RECT  2.350 1.010 4.035 1.100 ;
        RECT  2.250 0.500 2.350 1.100 ;
        RECT  0.950 0.500 2.250 0.590 ;
        RECT  0.950 1.210 1.005 1.300 ;
        RECT  0.045 0.500 0.450 0.590 ;
        RECT  0.295 1.210 0.450 1.300 ;
        RECT  4.820 1.030 4.925 1.490 ;
        RECT  3.880 1.390 4.820 1.490 ;
        RECT  2.545 0.500 4.705 0.590 ;
        RECT  3.780 1.210 3.880 1.490 ;
        RECT  2.665 1.210 3.780 1.300 ;
        RECT  2.455 0.310 2.545 0.590 ;
        RECT  0.295 0.310 2.455 0.410 ;
        RECT  1.225 1.210 2.335 1.300 ;
        RECT  1.120 1.030 1.225 1.490 ;
        RECT  0.180 1.390 1.120 1.490 ;
        RECT  0.060 1.240 0.180 1.490 ;
    END
END OAI22D4

MACRO OAI31D0
    CLASS CORE ;
    FOREIGN OAI31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.350 1.300 ;
        RECT  0.185 0.510 1.250 0.605 ;
        RECT  0.945 1.210 1.250 1.300 ;
        RECT  0.835 1.210 0.945 1.490 ;
        RECT  0.050 0.280 0.185 0.605 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.930 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.790 0.930 ;
        RECT  0.650 0.710 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.165 1.400 0.165 ;
        RECT  1.150 -0.165 1.320 0.405 ;
        RECT  0.000 -0.165 1.150 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.635 1.400 1.965 ;
        RECT  1.090 1.410 1.260 1.965 ;
        RECT  0.200 1.635 1.090 1.965 ;
        RECT  0.080 1.335 0.200 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.285 0.310 1.045 0.420 ;
    END
END OAI31D0

MACRO OAI31D1
    CLASS CORE ;
    FOREIGN OAI31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.500 1.350 1.300 ;
        RECT  0.045 0.500 1.250 0.590 ;
        RECT  0.795 1.210 1.250 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.950 0.700 1.050 0.950 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.165 1.400 0.165 ;
        RECT  1.110 -0.165 1.280 0.390 ;
        RECT  0.000 -0.165 1.110 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.635 1.400 1.965 ;
        RECT  1.090 1.410 1.260 1.965 ;
        RECT  0.200 1.635 1.090 1.965 ;
        RECT  0.080 1.335 0.200 1.965 ;
        RECT  0.000 1.635 0.080 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.285 0.310 1.000 0.410 ;
    END
END OAI31D1

MACRO OAI31D2
    CLASS CORE ;
    FOREIGN OAI31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4420 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.570 2.350 1.300 ;
        RECT  1.555 0.570 2.250 0.660 ;
        RECT  1.530 1.210 2.250 1.300 ;
        RECT  1.450 0.500 1.555 0.660 ;
        RECT  1.440 1.210 1.530 1.490 ;
        RECT  0.300 0.500 1.450 0.590 ;
        RECT  0.805 1.390 1.440 1.490 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.900 2.150 1.100 ;
        RECT  1.850 0.760 1.950 1.100 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.700 0.950 0.900 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.700 1.350 0.900 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.550 1.010 1.050 1.100 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.760 1.620 0.960 ;
        RECT  1.450 0.760 1.550 1.100 ;
        RECT  1.330 1.010 1.450 1.100 ;
        RECT  1.240 1.010 1.330 1.300 ;
        RECT  0.360 1.210 1.240 1.300 ;
        RECT  0.270 1.020 0.360 1.300 ;
        RECT  0.170 1.020 0.270 1.120 ;
        RECT  0.050 0.680 0.170 1.120 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.080 -0.165 2.400 0.165 ;
        RECT  1.900 -0.165 2.080 0.300 ;
        RECT  0.000 -0.165 1.900 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.635 2.400 1.965 ;
        RECT  1.640 1.390 1.820 1.965 ;
        RECT  0.175 1.635 1.640 1.965 ;
        RECT  0.055 1.230 0.175 1.965 ;
        RECT  0.000 1.635 0.055 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.220 0.285 2.340 0.480 ;
        RECT  1.790 0.390 2.220 0.480 ;
        RECT  1.650 0.310 1.790 0.480 ;
        RECT  0.190 0.310 1.650 0.410 ;
        RECT  0.085 0.310 0.190 0.560 ;
    END
END OAI31D2

MACRO OAI31D4
    CLASS CORE ;
    FOREIGN OAI31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.210 4.460 1.300 ;
        RECT  3.650 0.950 3.750 1.300 ;
        RECT  3.350 0.950 3.650 1.050 ;
        RECT  3.350 0.500 3.390 0.590 ;
        RECT  3.250 0.500 3.350 1.050 ;
        RECT  1.050 0.500 3.250 0.590 ;
        RECT  0.750 0.500 1.050 1.300 ;
        RECT  0.070 0.500 0.750 0.590 ;
        RECT  0.340 1.210 0.750 1.300 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.995 0.710 4.405 0.890 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.710 0.605 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.595 0.710 2.005 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.710 3.005 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.170 -0.165 4.800 0.165 ;
        RECT  4.170 0.310 4.460 0.410 ;
        RECT  4.030 -0.165 4.170 0.410 ;
        RECT  0.000 -0.165 4.030 0.165 ;
        RECT  3.750 0.310 4.030 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.635 4.800 1.965 ;
        RECT  4.570 1.030 4.680 1.965 ;
        RECT  3.370 1.635 4.570 1.965 ;
        RECT  3.370 1.390 4.210 1.500 ;
        RECT  3.220 1.390 3.370 1.965 ;
        RECT  2.460 1.390 3.220 1.500 ;
        RECT  0.000 1.635 3.220 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.750 1.210 4.460 1.300 ;
        RECT  3.650 0.950 3.750 1.300 ;
        RECT  3.350 0.950 3.650 1.050 ;
        RECT  3.350 0.500 3.390 0.590 ;
        RECT  3.250 0.500 3.350 1.050 ;
        RECT  1.150 0.500 3.250 0.590 ;
        RECT  0.070 0.500 0.650 0.590 ;
        RECT  0.340 1.210 0.650 1.300 ;
        RECT  4.575 0.350 4.680 0.590 ;
        RECT  3.635 0.500 4.575 0.590 ;
        RECT  3.535 0.310 3.635 0.590 ;
        RECT  0.330 0.310 3.535 0.410 ;
        RECT  1.370 1.210 3.420 1.300 ;
        RECT  0.225 1.390 2.340 1.500 ;
        RECT  0.120 1.150 0.225 1.500 ;
    END
END OAI31D4

MACRO OAI32D0
    CLASS CORE ;
    FOREIGN OAI32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 1.210 0.985 1.505 ;
        RECT  0.150 1.210 0.835 1.300 ;
        RECT  0.190 0.500 0.775 0.600 ;
        RECT  0.150 0.280 0.190 0.600 ;
        RECT  0.050 0.280 0.150 1.300 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.150 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.700 1.395 0.910 ;
        RECT  1.250 0.700 1.350 1.100 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.950 1.100 ;
        RECT  0.745 0.710 0.850 0.930 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.580 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.710 0.350 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 1.600 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.635 1.600 1.965 ;
        RECT  1.380 1.295 1.490 1.965 ;
        RECT  0.170 1.635 1.380 1.965 ;
        RECT  0.170 1.410 0.250 1.520 ;
        RECT  0.060 1.410 0.170 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.300 1.550 0.410 ;
    END
END OAI32D0

MACRO OAI32D1
    CLASS CORE ;
    FOREIGN OAI32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.210 0.995 1.490 ;
        RECT  0.150 1.210 0.830 1.300 ;
        RECT  0.150 0.500 0.750 0.590 ;
        RECT  0.050 0.500 0.150 1.300 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.700 1.150 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.700 1.395 0.910 ;
        RECT  1.250 0.700 1.350 1.100 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.700 0.950 1.100 ;
        RECT  0.740 0.700 0.850 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.580 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.700 0.350 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.165 1.600 0.165 ;
        RECT  1.080 -0.165 1.270 0.410 ;
        RECT  0.000 -0.165 1.080 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.495 1.635 1.600 1.965 ;
        RECT  1.375 1.210 1.495 1.965 ;
        RECT  0.220 1.635 1.375 1.965 ;
        RECT  0.050 1.410 0.220 1.965 ;
        RECT  0.000 1.635 0.050 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.965 0.500 1.530 0.590 ;
        RECT  0.865 0.310 0.965 0.590 ;
        RECT  0.300 0.310 0.865 0.410 ;
    END
END OAI32D1

MACRO OAI32D2
    CLASS CORE ;
    FOREIGN OAI32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4420 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.505 2.950 1.495 ;
        RECT  1.360 0.505 2.850 0.600 ;
        RECT  0.750 1.395 2.850 1.495 ;
        RECT  0.625 1.200 0.750 1.495 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.750 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.780 1.140 0.890 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.350 1.000 0.850 1.090 ;
        RECT  0.250 0.710 0.350 1.090 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.710 2.150 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.375 1.090 ;
        RECT  1.750 1.000 2.250 1.090 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.450 0.710 1.650 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.730 2.655 1.290 ;
        RECT  1.350 1.200 2.545 1.290 ;
        RECT  1.250 0.710 1.350 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.165 3.000 0.165 ;
        RECT  0.770 0.295 1.050 0.400 ;
        RECT  0.630 -0.165 0.770 0.400 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.315 0.295 0.630 0.400 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.215 1.635 3.000 1.965 ;
        RECT  0.105 1.200 0.215 1.965 ;
        RECT  0.000 1.635 0.105 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.295 2.880 0.395 ;
        RECT  1.160 0.295 1.250 0.600 ;
        RECT  0.060 0.500 1.160 0.600 ;
    END
END OAI32D2

MACRO OAI32D4
    CLASS CORE ;
    FOREIGN OAI32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.510 2.915 0.620 ;
        RECT  2.850 1.110 2.915 1.220 ;
        RECT  2.550 0.510 2.850 1.220 ;
        RECT  2.185 0.510 2.550 0.620 ;
        RECT  2.185 1.110 2.550 1.220 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.160 1.090 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.710 1.405 0.940 ;
        RECT  1.250 0.710 1.350 1.090 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.710 0.950 1.090 ;
        RECT  0.775 0.710 0.850 0.940 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.565 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.125 -0.165 3.200 0.165 ;
        RECT  3.015 -0.165 3.125 0.695 ;
        RECT  2.370 -0.165 3.015 0.165 ;
        RECT  2.370 0.305 2.655 0.415 ;
        RECT  2.230 -0.165 2.370 0.415 ;
        RECT  1.290 -0.165 2.230 0.165 ;
        RECT  1.925 0.305 2.230 0.415 ;
        RECT  1.080 -0.165 1.290 0.410 ;
        RECT  0.000 -0.165 1.080 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.125 1.635 3.200 1.965 ;
        RECT  3.015 1.040 3.125 1.965 ;
        RECT  2.370 1.635 3.015 1.965 ;
        RECT  2.370 1.330 2.655 1.440 ;
        RECT  2.230 1.330 2.370 1.965 ;
        RECT  1.925 1.330 2.230 1.440 ;
        RECT  0.970 1.635 2.230 1.965 ;
        RECT  0.970 1.390 1.550 1.495 ;
        RECT  0.830 1.390 0.970 1.965 ;
        RECT  0.050 1.390 0.830 1.495 ;
        RECT  0.000 1.635 0.830 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.185 0.510 2.450 0.620 ;
        RECT  2.185 1.110 2.450 1.220 ;
        RECT  2.075 0.775 2.340 0.890 ;
        RECT  1.985 0.585 2.075 1.150 ;
        RECT  1.825 0.585 1.985 0.695 ;
        RECT  1.825 1.040 1.985 1.150 ;
        RECT  1.605 0.785 1.875 0.890 ;
        RECT  1.715 0.295 1.825 0.695 ;
        RECT  1.715 1.040 1.825 1.470 ;
        RECT  1.515 0.785 1.605 1.300 ;
        RECT  0.970 0.500 1.550 0.600 ;
        RECT  0.360 1.200 1.515 1.300 ;
        RECT  0.880 0.310 0.970 0.600 ;
        RECT  0.300 0.310 0.880 0.410 ;
        RECT  0.360 0.500 0.770 0.600 ;
        RECT  0.270 0.500 0.360 1.300 ;
        RECT  0.060 0.500 0.270 0.600 ;
    END
END OAI32D4

MACRO OAI32XD4
    CLASS CORE ;
    FOREIGN OAI32XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.500 5.495 0.600 ;
        RECT  3.850 1.000 5.485 1.115 ;
        RECT  3.550 0.500 3.850 1.115 ;
        RECT  2.425 0.500 3.550 0.600 ;
        RECT  3.320 1.000 3.550 1.115 ;
        RECT  3.210 1.000 3.320 1.305 ;
        RECT  0.605 1.205 3.210 1.305 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.710 1.950 0.890 ;
        RECT  1.650 0.710 1.760 1.115 ;
        RECT  0.950 1.000 1.650 1.115 ;
        RECT  0.840 0.710 0.950 1.115 ;
        RECT  0.650 0.710 0.840 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2201 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.500 2.160 0.940 ;
        RECT  1.355 0.500 2.050 0.600 ;
        RECT  1.245 0.500 1.355 0.910 ;
        RECT  0.350 0.500 1.245 0.600 ;
        RECT  0.240 0.500 0.350 0.940 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.710 5.205 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.995 0.710 4.405 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2191 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.710 3.005 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 5.800 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.635 5.800 1.965 ;
        RECT  1.770 1.395 2.355 1.505 ;
        RECT  1.630 1.395 1.770 1.965 ;
        RECT  1.125 1.395 1.630 1.505 ;
        RECT  0.245 1.635 1.630 1.965 ;
        RECT  0.135 1.040 0.245 1.965 ;
        RECT  0.000 1.635 0.135 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.950 0.500 5.495 0.600 ;
        RECT  3.950 1.000 5.485 1.115 ;
        RECT  2.425 0.500 3.450 0.600 ;
        RECT  3.320 1.000 3.450 1.115 ;
        RECT  3.210 1.000 3.320 1.305 ;
        RECT  0.605 1.205 3.210 1.305 ;
        RECT  0.085 0.300 5.745 0.410 ;
        RECT  5.595 1.040 5.705 1.470 ;
        RECT  3.465 1.205 5.595 1.305 ;
        RECT  2.445 1.395 4.455 1.505 ;
    END
END OAI32XD4

MACRO OAI33D0
    CLASS CORE ;
    FOREIGN OAI33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 1.310 1.010 1.490 ;
        RECT  0.350 0.495 0.755 0.600 ;
        RECT  0.450 1.210 0.545 1.490 ;
        RECT  0.350 1.210 0.450 1.300 ;
        RECT  0.260 0.495 0.350 1.300 ;
        RECT  0.180 0.495 0.260 0.590 ;
        RECT  0.050 0.280 0.180 0.590 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.090 ;
        RECT  1.030 0.700 1.050 0.910 ;
        RECT  0.940 0.740 1.030 0.910 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.680 1.350 1.110 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.910 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0354 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.790 0.950 ;
        RECT  0.650 0.710 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0354 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.490 ;
        RECT  0.000 -0.165 1.615 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.635 1.800 1.965 ;
        RECT  1.605 1.300 1.715 1.965 ;
        RECT  0.340 1.635 1.605 1.965 ;
        RECT  0.240 1.390 0.340 1.965 ;
        RECT  0.050 1.390 0.240 1.495 ;
        RECT  0.000 1.635 0.240 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.285 0.295 1.515 0.405 ;
    END
END OAI33D0

MACRO OAI33D1
    CLASS CORE ;
    FOREIGN OAI33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 1.310 1.010 1.490 ;
        RECT  0.350 0.500 0.755 0.590 ;
        RECT  0.450 1.210 0.545 1.490 ;
        RECT  0.350 1.210 0.450 1.300 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 0.500 0.260 0.590 ;
        RECT  0.075 0.310 0.180 0.590 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.090 ;
        RECT  1.030 0.700 1.050 0.910 ;
        RECT  0.940 0.740 1.030 0.910 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.680 1.350 1.110 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.910 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.165 1.800 0.165 ;
        RECT  1.615 -0.165 1.725 0.565 ;
        RECT  0.000 -0.165 1.615 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.635 1.800 1.965 ;
        RECT  1.605 1.070 1.715 1.965 ;
        RECT  0.340 1.635 1.605 1.965 ;
        RECT  0.240 1.390 0.340 1.965 ;
        RECT  0.050 1.390 0.240 1.495 ;
        RECT  0.000 1.635 0.240 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.295 0.310 1.500 0.410 ;
    END
END OAI33D1

MACRO OAI33D2
    CLASS CORE ;
    FOREIGN OAI33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4420 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.510 3.350 1.490 ;
        RECT  1.810 0.510 3.250 0.600 ;
        RECT  0.800 1.390 3.250 1.490 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.700 0.950 0.900 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1104 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.700 1.350 0.900 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.550 1.010 1.050 1.100 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.710 1.560 1.100 ;
        RECT  1.365 1.010 1.440 1.100 ;
        RECT  1.260 1.010 1.365 1.300 ;
        RECT  0.360 1.210 1.260 1.300 ;
        RECT  0.270 1.020 0.360 1.300 ;
        RECT  0.170 1.020 0.270 1.120 ;
        RECT  0.050 0.680 0.170 1.120 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.550 0.900 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.825 1.100 ;
        RECT  2.150 1.010 2.650 1.100 ;
        RECT  1.985 0.710 2.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.020 0.710 3.155 1.290 ;
        RECT  1.805 1.190 3.020 1.290 ;
        RECT  1.650 0.710 1.805 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.165 3.400 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 1.635 3.400 1.965 ;
        RECT  0.060 1.230 0.180 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.700 0.300 3.300 0.400 ;
        RECT  1.590 0.300 1.700 0.520 ;
        RECT  0.050 0.410 1.590 0.520 ;
    END
END OAI33D2

MACRO OAI33D4
    CLASS CORE ;
    FOREIGN OAI33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.310 2.645 0.420 ;
        RECT  2.450 0.995 2.630 1.115 ;
        RECT  2.150 0.310 2.450 1.115 ;
        RECT  1.900 0.310 2.150 0.420 ;
        RECT  1.900 0.995 2.150 1.115 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.100 ;
        RECT  0.940 0.700 1.050 0.910 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.700 1.380 1.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.700 1.755 1.100 ;
        RECT  1.530 0.700 1.645 0.910 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.700 0.790 0.950 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.865 -0.165 3.200 0.165 ;
        RECT  2.755 -0.165 2.865 0.455 ;
        RECT  1.780 -0.165 2.755 0.165 ;
        RECT  1.630 -0.165 1.780 0.580 ;
        RECT  0.000 -0.165 1.630 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.635 3.200 1.965 ;
        RECT  2.370 1.390 2.905 1.490 ;
        RECT  2.230 1.390 2.370 1.965 ;
        RECT  1.585 1.390 2.230 1.490 ;
        RECT  0.330 1.635 2.230 1.965 ;
        RECT  0.230 1.390 0.330 1.965 ;
        RECT  0.055 1.390 0.230 1.495 ;
        RECT  0.000 1.635 0.230 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.310 2.645 0.420 ;
        RECT  2.550 0.995 2.630 1.115 ;
        RECT  1.900 0.310 2.050 0.420 ;
        RECT  1.900 0.995 2.050 1.115 ;
        RECT  3.060 0.280 3.150 1.490 ;
        RECT  3.015 0.280 3.060 0.655 ;
        RECT  3.015 1.040 3.060 1.490 ;
        RECT  2.695 0.565 3.015 0.655 ;
        RECT  2.900 0.765 2.950 0.935 ;
        RECT  2.810 0.765 2.900 1.300 ;
        RECT  0.975 1.210 2.810 1.300 ;
        RECT  2.585 0.565 2.695 0.895 ;
        RECT  0.290 0.310 1.515 0.410 ;
        RECT  0.825 1.210 0.975 1.420 ;
        RECT  0.350 1.210 0.825 1.300 ;
        RECT  0.350 0.500 0.755 0.590 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.180 0.500 0.260 0.590 ;
        RECT  0.075 0.350 0.180 0.590 ;
    END
END OAI33D4

MACRO OAI33XD4
    CLASS CORE ;
    FOREIGN OAI33XD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.500 6.715 0.600 ;
        RECT  5.250 1.000 6.715 1.115 ;
        RECT  4.950 0.500 5.250 1.115 ;
        RECT  3.645 0.500 4.950 0.600 ;
        RECT  0.285 1.000 4.950 1.115 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.950 0.890 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.950 0.890 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2186 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 3.150 0.890 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.710 6.550 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.710 5.750 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.165 7.000 0.165 ;
        RECT  2.970 0.300 3.315 0.410 ;
        RECT  2.830 -0.165 2.970 0.410 ;
        RECT  1.770 -0.165 2.830 0.165 ;
        RECT  2.615 0.300 2.830 0.410 ;
        RECT  1.770 0.300 2.045 0.410 ;
        RECT  1.630 -0.165 1.770 0.410 ;
        RECT  0.770 -0.165 1.630 0.165 ;
        RECT  1.335 0.300 1.630 0.410 ;
        RECT  0.770 0.300 1.005 0.410 ;
        RECT  0.630 -0.165 0.770 0.410 ;
        RECT  0.000 -0.165 0.630 0.165 ;
        RECT  0.295 0.300 0.630 0.410 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.370 1.635 7.000 1.965 ;
        RECT  4.370 1.395 4.615 1.505 ;
        RECT  4.230 1.395 4.370 1.965 ;
        RECT  3.905 1.395 4.230 1.505 ;
        RECT  3.370 1.635 4.230 1.965 ;
        RECT  3.370 1.395 3.595 1.505 ;
        RECT  3.230 1.395 3.370 1.965 ;
        RECT  2.865 1.395 3.230 1.505 ;
        RECT  0.000 1.635 3.230 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.350 0.500 6.715 0.600 ;
        RECT  5.350 1.000 6.715 1.115 ;
        RECT  3.645 0.500 4.850 0.600 ;
        RECT  0.285 1.000 4.850 1.115 ;
        RECT  6.825 0.300 6.935 0.510 ;
        RECT  6.815 1.040 6.925 1.505 ;
        RECT  3.535 0.300 6.825 0.410 ;
        RECT  4.705 1.395 6.815 1.505 ;
        RECT  3.655 1.205 5.675 1.305 ;
        RECT  3.425 0.300 3.535 0.600 ;
        RECT  2.505 0.500 3.425 0.600 ;
        RECT  1.325 1.205 3.325 1.305 ;
        RECT  2.395 0.275 2.505 0.695 ;
        RECT  2.265 0.500 2.395 0.600 ;
        RECT  0.185 1.395 2.315 1.505 ;
        RECT  2.155 0.275 2.265 0.695 ;
        RECT  1.225 0.500 2.155 0.600 ;
        RECT  1.115 0.275 1.225 0.695 ;
        RECT  0.185 0.500 1.115 0.600 ;
        RECT  0.075 0.275 0.185 0.695 ;
        RECT  0.075 1.040 0.185 1.505 ;
    END
END OAI33XD4

MACRO OD18DCAP16
    CLASS CORE ;
    FOREIGN OD18DCAP16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.535 -0.165 3.200 0.165 ;
        RECT  2.385 -0.165 2.535 1.145 ;
        RECT  0.815 -0.165 2.385 0.165 ;
        RECT  0.665 -0.165 0.815 1.145 ;
        RECT  0.000 -0.165 0.665 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.595 1.635 3.200 1.965 ;
        RECT  1.595 1.305 2.305 1.455 ;
        RECT  1.405 1.305 1.595 1.965 ;
        RECT  0.895 1.305 1.405 1.455 ;
        RECT  0.000 1.635 1.405 1.965 ;
        END
    END VDD
END OD18DCAP16

MACRO OD18DCAP32
    CLASS CORE ;
    FOREIGN OD18DCAP32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.735 -0.165 6.400 0.165 ;
        RECT  5.585 -0.165 5.735 1.145 ;
        RECT  3.285 -0.165 5.585 0.165 ;
        RECT  3.115 -0.165 3.285 1.145 ;
        RECT  0.810 -0.165 3.115 0.165 ;
        RECT  0.665 -0.165 0.810 1.145 ;
        RECT  0.000 -0.165 0.665 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.595 1.635 6.400 1.965 ;
        RECT  4.595 1.305 5.505 1.455 ;
        RECT  4.405 1.305 4.595 1.965 ;
        RECT  3.355 1.305 4.405 1.455 ;
        RECT  1.995 1.635 4.405 1.965 ;
        RECT  1.995 1.305 3.045 1.455 ;
        RECT  1.805 1.305 1.995 1.965 ;
        RECT  0.895 1.305 1.805 1.455 ;
        RECT  0.000 1.635 1.805 1.965 ;
        END
    END VDD
END OD18DCAP32

MACRO OD18DCAP64
    CLASS CORE ;
    FOREIGN OD18DCAP64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.135 -0.165 12.800 0.165 ;
        RECT  11.985 -0.165 12.135 1.145 ;
        RECT  9.325 -0.165 11.985 0.165 ;
        RECT  9.135 -0.165 9.325 1.145 ;
        RECT  6.485 -0.165 9.135 0.165 ;
        RECT  6.315 -0.165 6.485 1.145 ;
        RECT  3.665 -0.165 6.315 0.165 ;
        RECT  3.475 -0.165 3.665 1.145 ;
        RECT  0.805 -0.165 3.475 0.165 ;
        RECT  0.645 -0.165 0.805 1.145 ;
        RECT  0.000 -0.165 0.645 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.795 1.635 12.800 1.965 ;
        RECT  10.795 1.305 11.905 1.455 ;
        RECT  10.605 1.305 10.795 1.965 ;
        RECT  9.385 1.305 10.605 1.455 ;
        RECT  7.995 1.635 10.605 1.965 ;
        RECT  7.995 1.305 9.075 1.455 ;
        RECT  7.805 1.305 7.995 1.965 ;
        RECT  6.555 1.305 7.805 1.455 ;
        RECT  5.195 1.635 7.805 1.965 ;
        RECT  5.195 1.305 6.245 1.455 ;
        RECT  5.005 1.305 5.195 1.965 ;
        RECT  3.725 1.305 5.005 1.455 ;
        RECT  2.195 1.635 5.005 1.965 ;
        RECT  2.195 1.305 3.415 1.455 ;
        RECT  2.005 1.305 2.195 1.965 ;
        RECT  0.895 1.305 2.005 1.455 ;
        RECT  0.000 1.635 2.005 1.965 ;
        END
    END VDD
END OD18DCAP64

MACRO OR2D0
    CLASS CORE ;
    FOREIGN OR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.485 1.150 1.500 ;
        RECT  0.995 0.485 1.050 0.685 ;
        RECT  0.995 1.300 1.050 1.500 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.780 0.660 0.890 ;
        RECT  0.450 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.755 0.350 0.920 ;
        RECT  0.050 0.500 0.150 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 -0.165 1.200 0.165 ;
        RECT  0.680 -0.165 0.850 0.390 ;
        RECT  0.270 -0.165 0.680 0.165 ;
        RECT  0.100 -0.165 0.270 0.390 ;
        RECT  0.000 -0.165 0.100 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.635 1.200 1.965 ;
        RECT  0.660 1.410 0.830 1.965 ;
        RECT  0.000 1.635 0.660 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 0.780 0.940 0.890 ;
        RECT  0.770 0.500 0.860 1.320 ;
        RECT  0.370 0.500 0.770 0.600 ;
        RECT  0.245 1.210 0.770 1.320 ;
        RECT  0.135 1.210 0.245 1.470 ;
    END
END OR2D0

MACRO OR2D1
    CLASS CORE ;
    FOREIGN OR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.300 1.150 1.500 ;
        RECT  0.995 0.300 1.050 0.685 ;
        RECT  0.995 1.100 1.050 1.500 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0437 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.780 0.660 0.890 ;
        RECT  0.450 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0434 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.755 0.350 0.920 ;
        RECT  0.050 0.500 0.150 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 -0.165 1.200 0.165 ;
        RECT  0.680 -0.165 0.850 0.390 ;
        RECT  0.270 -0.165 0.680 0.165 ;
        RECT  0.100 -0.165 0.270 0.390 ;
        RECT  0.000 -0.165 0.100 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.635 1.200 1.965 ;
        RECT  0.660 1.410 0.830 1.965 ;
        RECT  0.000 1.635 0.660 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 0.780 0.940 0.890 ;
        RECT  0.770 0.500 0.860 1.320 ;
        RECT  0.370 0.500 0.770 0.600 ;
        RECT  0.245 1.210 0.770 1.320 ;
        RECT  0.135 1.040 0.245 1.470 ;
    END
END OR2D1

MACRO OR2D2
    CLASS CORE ;
    FOREIGN OR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.575 1.150 1.170 ;
        RECT  0.940 0.295 1.050 0.685 ;
        RECT  1.040 1.060 1.050 1.170 ;
        RECT  0.930 1.060 1.040 1.470 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0437 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.700 0.605 0.920 ;
        RECT  0.450 0.700 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.240 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 -0.165 1.400 0.165 ;
        RECT  1.195 -0.165 1.315 0.475 ;
        RECT  0.795 -0.165 1.195 0.165 ;
        RECT  0.625 -0.165 0.795 0.390 ;
        RECT  0.190 -0.165 0.625 0.165 ;
        RECT  0.070 -0.165 0.190 0.590 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 1.635 1.400 1.965 ;
        RECT  1.195 1.325 1.315 1.965 ;
        RECT  0.775 1.635 1.195 1.965 ;
        RECT  0.605 1.410 0.775 1.965 ;
        RECT  0.000 1.635 0.605 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.840 0.750 0.875 0.920 ;
        RECT  0.730 0.500 0.840 1.320 ;
        RECT  0.315 0.500 0.730 0.610 ;
        RECT  0.190 1.210 0.730 1.320 ;
        RECT  0.080 1.210 0.190 1.485 ;
    END
END OR2D2

MACRO OR2D4
    CLASS CORE ;
    FOREIGN OR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.035 0.275 2.065 0.695 ;
        RECT  2.035 1.040 2.065 1.490 ;
        RECT  1.955 0.275 2.035 1.490 ;
        RECT  1.750 0.545 1.955 1.190 ;
        RECT  1.540 0.545 1.750 0.695 ;
        RECT  1.540 1.040 1.750 1.190 ;
        RECT  1.440 0.275 1.540 0.695 ;
        RECT  1.430 1.040 1.540 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0869 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.150 1.500 ;
        RECT  0.485 1.410 1.040 1.500 ;
        RECT  0.385 1.000 0.485 1.500 ;
        RECT  0.350 1.000 0.385 1.100 ;
        RECT  0.250 0.700 0.350 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0858 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 -0.165 2.400 0.165 ;
        RECT  2.215 -0.165 2.325 0.695 ;
        RECT  1.805 -0.165 2.215 0.165 ;
        RECT  1.695 -0.165 1.805 0.455 ;
        RECT  0.785 -0.165 1.695 0.165 ;
        RECT  0.610 -0.165 0.785 0.410 ;
        RECT  0.210 -0.165 0.610 0.165 ;
        RECT  0.100 -0.165 0.210 0.475 ;
        RECT  0.000 -0.165 0.100 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 1.635 2.400 1.965 ;
        RECT  2.215 1.040 2.325 1.965 ;
        RECT  1.800 1.635 2.215 1.965 ;
        RECT  1.690 1.280 1.800 1.965 ;
        RECT  0.230 1.635 1.690 1.965 ;
        RECT  0.120 1.210 0.230 1.965 ;
        RECT  0.000 1.635 0.120 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.540 0.545 1.650 0.695 ;
        RECT  1.540 1.040 1.650 1.190 ;
        RECT  1.440 0.275 1.540 0.695 ;
        RECT  1.430 1.040 1.540 1.490 ;
        RECT  1.330 0.785 1.535 0.890 ;
        RECT  1.240 0.500 1.330 0.890 ;
        RECT  1.035 0.500 1.240 0.590 ;
        RECT  0.930 0.275 1.035 0.590 ;
        RECT  0.920 0.275 0.930 1.320 ;
        RECT  0.840 0.500 0.920 1.320 ;
        RECT  0.470 0.500 0.840 0.590 ;
        RECT  0.595 1.210 0.840 1.320 ;
        RECT  0.360 0.275 0.470 0.590 ;
    END
END OR2D4

MACRO OR2D8
    CLASS CORE ;
    FOREIGN OR2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.295 3.465 0.690 ;
        RECT  3.350 1.050 3.465 1.490 ;
        RECT  2.955 0.585 3.350 0.690 ;
        RECT  2.955 1.050 3.350 1.160 ;
        RECT  2.845 0.295 2.955 0.690 ;
        RECT  2.845 1.050 2.955 1.460 ;
        RECT  2.650 0.585 2.845 0.690 ;
        RECT  2.650 1.050 2.845 1.160 ;
        RECT  2.455 0.585 2.650 1.160 ;
        RECT  2.350 0.295 2.455 1.460 ;
        RECT  2.345 0.295 2.350 0.690 ;
        RECT  2.345 1.050 2.350 1.460 ;
        RECT  1.955 0.585 2.345 0.690 ;
        RECT  1.955 1.050 2.345 1.160 ;
        RECT  1.845 0.295 1.955 0.690 ;
        RECT  1.845 1.050 1.955 1.460 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.1311 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.700 1.555 1.130 ;
        RECT  0.750 1.030 1.435 1.130 ;
        RECT  0.650 0.780 0.750 1.130 ;
        RECT  0.560 0.780 0.650 0.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1295 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.600 1.150 0.920 ;
        RECT  0.170 0.600 1.040 0.690 ;
        RECT  0.050 0.600 0.170 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.165 3.800 0.165 ;
        RECT  3.615 -0.165 3.725 0.685 ;
        RECT  0.190 -0.165 3.615 0.165 ;
        RECT  0.070 -0.165 0.190 0.475 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 1.635 3.800 1.965 ;
        RECT  3.615 1.050 3.725 1.965 ;
        RECT  0.000 1.635 3.615 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.350 0.295 3.465 0.690 ;
        RECT  3.350 1.050 3.465 1.490 ;
        RECT  2.955 0.585 3.350 0.690 ;
        RECT  2.955 1.050 3.350 1.160 ;
        RECT  2.845 0.295 2.955 0.690 ;
        RECT  2.845 1.050 2.955 1.460 ;
        RECT  2.750 0.585 2.845 0.690 ;
        RECT  2.750 1.050 2.845 1.160 ;
        RECT  1.955 0.585 2.250 0.690 ;
        RECT  1.955 1.050 2.250 1.160 ;
        RECT  1.845 0.295 1.955 0.690 ;
        RECT  1.845 1.050 1.955 1.460 ;
        RECT  2.830 0.780 3.475 0.890 ;
        RECT  1.745 0.780 2.170 0.890 ;
        RECT  1.645 0.420 1.745 1.350 ;
        RECT  1.475 0.420 1.645 0.510 ;
        RECT  0.185 1.240 1.645 1.350 ;
        RECT  1.325 0.275 1.475 0.510 ;
        RECT  0.965 0.420 1.325 0.510 ;
        RECT  0.815 0.275 0.965 0.510 ;
        RECT  0.465 0.420 0.815 0.510 ;
        RECT  0.315 0.275 0.465 0.510 ;
        RECT  0.075 1.240 0.185 1.470 ;
    END
END OR2D8

MACRO OR2XD1
    CLASS CORE ;
    FOREIGN OR2XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.300 1.150 1.500 ;
        RECT  0.995 0.300 1.050 0.685 ;
        RECT  0.995 1.100 1.050 1.500 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.780 0.660 0.890 ;
        RECT  0.450 0.710 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.755 0.350 0.920 ;
        RECT  0.050 0.500 0.150 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 -0.165 1.200 0.165 ;
        RECT  0.680 -0.165 0.850 0.390 ;
        RECT  0.270 -0.165 0.680 0.165 ;
        RECT  0.100 -0.165 0.270 0.390 ;
        RECT  0.000 -0.165 0.100 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.635 1.200 1.965 ;
        RECT  0.660 1.410 0.830 1.965 ;
        RECT  0.000 1.635 0.660 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 0.780 0.940 0.890 ;
        RECT  0.770 0.500 0.860 1.320 ;
        RECT  0.370 0.500 0.770 0.600 ;
        RECT  0.245 1.210 0.770 1.320 ;
        RECT  0.135 1.040 0.245 1.470 ;
    END
END OR2XD1

MACRO OR3D0
    CLASS CORE ;
    FOREIGN OR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.295 1.350 1.490 ;
        RECT  1.215 0.295 1.250 0.485 ;
        RECT  1.195 1.260 1.250 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.350 1.100 ;
        RECT  0.150 0.780 0.250 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.750 0.850 0.920 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.165 1.400 0.165 ;
        RECT  0.900 -0.165 1.070 0.410 ;
        RECT  0.500 -0.165 0.900 0.165 ;
        RECT  0.330 -0.165 0.500 0.410 ;
        RECT  0.000 -0.165 0.330 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.635 1.400 1.965 ;
        RECT  0.880 1.410 1.050 1.965 ;
        RECT  0.000 1.635 0.880 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.035 0.750 1.130 0.920 ;
        RECT  0.945 0.500 1.035 1.320 ;
        RECT  0.755 0.500 0.945 0.590 ;
        RECT  0.205 1.210 0.945 1.320 ;
        RECT  0.645 0.295 0.755 0.590 ;
        RECT  0.185 0.500 0.645 0.590 ;
        RECT  0.095 1.210 0.205 1.490 ;
        RECT  0.075 0.305 0.185 0.590 ;
    END
END OR3D0

MACRO OR3D1
    CLASS CORE ;
    FOREIGN OR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.295 1.350 1.490 ;
        RECT  1.215 0.295 1.250 0.685 ;
        RECT  1.195 1.050 1.250 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.350 1.100 ;
        RECT  0.150 0.780 0.250 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.750 0.850 0.920 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.165 1.400 0.165 ;
        RECT  0.900 -0.165 1.070 0.410 ;
        RECT  0.500 -0.165 0.900 0.165 ;
        RECT  0.330 -0.165 0.500 0.410 ;
        RECT  0.000 -0.165 0.330 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.635 1.400 1.965 ;
        RECT  0.880 1.410 1.050 1.965 ;
        RECT  0.000 1.635 0.880 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.035 0.750 1.130 0.920 ;
        RECT  0.945 0.500 1.035 1.320 ;
        RECT  0.755 0.500 0.945 0.590 ;
        RECT  0.065 1.210 0.945 1.320 ;
        RECT  0.645 0.295 0.755 0.590 ;
        RECT  0.185 0.500 0.645 0.590 ;
        RECT  0.075 0.305 0.185 0.590 ;
    END
END OR3D1

MACRO OR3D2
    CLASS CORE ;
    FOREIGN OR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.565 1.350 1.125 ;
        RECT  1.250 0.275 1.265 1.490 ;
        RECT  1.155 0.275 1.250 0.695 ;
        RECT  1.155 1.030 1.250 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.710 0.180 0.920 ;
        RECT  0.050 0.710 0.150 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.560 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0437 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.850 0.920 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 -0.165 1.600 0.165 ;
        RECT  1.415 -0.165 1.525 0.465 ;
        RECT  0.500 -0.165 1.415 0.165 ;
        RECT  0.330 -0.165 0.500 0.410 ;
        RECT  0.000 -0.165 0.330 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 1.635 1.600 1.965 ;
        RECT  1.415 1.270 1.525 1.965 ;
        RECT  0.925 1.635 1.415 1.965 ;
        RECT  0.925 1.390 1.045 1.495 ;
        RECT  0.835 1.390 0.925 1.965 ;
        RECT  0.000 1.635 0.835 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.785 1.140 0.890 ;
        RECT  0.960 0.500 1.050 1.300 ;
        RECT  0.770 0.500 0.960 0.590 ;
        RECT  0.065 1.200 0.960 1.300 ;
        RECT  0.630 0.295 0.770 0.590 ;
        RECT  0.185 0.500 0.630 0.590 ;
        RECT  0.075 0.295 0.185 0.590 ;
    END
END OR3D2

MACRO OR3D4
    CLASS CORE ;
    FOREIGN OR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.275 2.465 0.685 ;
        RECT  2.450 1.050 2.465 1.490 ;
        RECT  2.355 0.275 2.450 1.490 ;
        RECT  2.150 0.585 2.355 1.150 ;
        RECT  1.945 0.585 2.150 0.695 ;
        RECT  1.945 1.050 2.150 1.150 ;
        RECT  1.840 0.275 1.945 0.695 ;
        RECT  1.840 1.050 1.945 1.460 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0866 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 0.790 0.950 1.100 ;
        RECT  0.650 0.900 0.760 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0866 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.585 1.290 0.940 ;
        RECT  0.550 0.585 1.180 0.685 ;
        RECT  0.450 0.585 0.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0869 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.710 1.550 1.300 ;
        RECT  0.340 1.210 1.430 1.300 ;
        RECT  0.250 0.980 0.340 1.300 ;
        RECT  0.180 0.980 0.250 1.090 ;
        RECT  0.050 0.700 0.180 1.090 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.725 -0.165 2.800 0.165 ;
        RECT  2.615 -0.165 2.725 0.685 ;
        RECT  2.205 -0.165 2.615 0.165 ;
        RECT  2.095 -0.165 2.205 0.495 ;
        RECT  0.185 -0.165 2.095 0.165 ;
        RECT  0.075 -0.165 0.185 0.485 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.725 1.635 2.800 1.965 ;
        RECT  2.615 1.050 2.725 1.965 ;
        RECT  2.205 1.635 2.615 1.965 ;
        RECT  2.095 1.240 2.205 1.965 ;
        RECT  0.170 1.635 2.095 1.965 ;
        RECT  0.170 1.390 0.250 1.495 ;
        RECT  0.060 1.390 0.170 1.965 ;
        RECT  0.000 1.635 0.060 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.945 0.585 2.050 0.695 ;
        RECT  1.945 1.050 2.050 1.150 ;
        RECT  1.840 0.275 1.945 0.695 ;
        RECT  1.840 1.050 1.945 1.460 ;
        RECT  1.750 0.805 2.000 0.915 ;
        RECT  1.660 0.325 1.750 1.495 ;
        RECT  0.285 0.325 1.660 0.435 ;
        RECT  0.760 1.390 1.660 1.495 ;
    END
END OR3D4

MACRO OR3D8
    CLASS CORE ;
    FOREIGN OR3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.155 0.275 4.265 0.685 ;
        RECT  4.155 1.050 4.265 1.460 ;
        RECT  3.765 0.585 4.155 0.685 ;
        RECT  3.765 1.050 4.155 1.160 ;
        RECT  3.655 0.275 3.765 0.685 ;
        RECT  3.655 1.050 3.765 1.460 ;
        RECT  3.450 0.585 3.655 0.685 ;
        RECT  3.450 1.050 3.655 1.160 ;
        RECT  3.245 0.585 3.450 1.160 ;
        RECT  3.150 0.275 3.245 1.460 ;
        RECT  3.140 0.275 3.150 0.685 ;
        RECT  3.135 1.050 3.150 1.460 ;
        RECT  2.745 0.585 3.140 0.685 ;
        RECT  2.745 1.050 3.135 1.160 ;
        RECT  2.635 0.275 2.745 0.685 ;
        RECT  2.635 1.050 2.745 1.460 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.1311 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.700 1.960 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.700 1.360 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.700 0.560 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 -0.165 4.600 0.165 ;
        RECT  4.415 -0.165 4.525 0.685 ;
        RECT  3.505 -0.165 4.415 0.165 ;
        RECT  3.395 -0.165 3.505 0.495 ;
        RECT  0.000 -0.165 3.395 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.635 4.600 1.965 ;
        RECT  4.415 1.050 4.525 1.965 ;
        RECT  3.505 1.635 4.415 1.965 ;
        RECT  3.395 1.250 3.505 1.965 ;
        RECT  0.000 1.635 3.395 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.155 0.275 4.265 0.685 ;
        RECT  4.155 1.050 4.265 1.460 ;
        RECT  3.765 0.585 4.155 0.685 ;
        RECT  3.765 1.050 4.155 1.160 ;
        RECT  3.655 0.275 3.765 0.685 ;
        RECT  3.655 1.050 3.765 1.460 ;
        RECT  3.550 0.585 3.655 0.685 ;
        RECT  3.550 1.050 3.655 1.160 ;
        RECT  2.635 0.275 2.745 0.685 ;
        RECT  2.635 1.050 2.745 1.460 ;
        RECT  2.295 0.780 3.030 0.890 ;
        RECT  2.190 0.325 2.295 0.890 ;
        RECT  2.135 1.050 2.245 1.460 ;
        RECT  0.800 0.325 2.190 0.435 ;
        RECT  1.745 1.190 2.135 1.300 ;
        RECT  1.635 1.050 1.745 1.460 ;
        RECT  1.065 1.190 1.635 1.300 ;
        RECT  0.295 1.390 1.525 1.495 ;
        RECT  0.700 0.325 0.800 1.300 ;
        RECT  0.045 0.325 0.700 0.435 ;
        RECT  0.185 1.190 0.700 1.300 ;
        RECT  0.075 1.050 0.185 1.460 ;
        RECT  2.745 0.585 3.050 0.685 ;
        RECT  2.745 1.050 3.050 1.160 ;
    END
END OR3D8

MACRO OR3XD1
    CLASS CORE ;
    FOREIGN OR3XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.295 1.350 1.490 ;
        RECT  1.215 0.295 1.250 0.685 ;
        RECT  1.195 1.050 1.250 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.700 0.350 1.100 ;
        RECT  0.150 0.780 0.250 0.890 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.700 0.560 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.750 0.850 0.920 ;
        RECT  0.650 0.700 0.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 -0.165 1.400 0.165 ;
        RECT  0.930 -0.165 1.040 0.410 ;
        RECT  0.470 -0.165 0.930 0.165 ;
        RECT  0.360 -0.165 0.470 0.410 ;
        RECT  0.000 -0.165 0.360 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.635 1.400 1.965 ;
        RECT  0.910 1.410 1.020 1.965 ;
        RECT  0.000 1.635 0.910 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.035 0.750 1.130 0.920 ;
        RECT  0.945 0.500 1.035 1.320 ;
        RECT  0.755 0.500 0.945 0.590 ;
        RECT  0.065 1.210 0.945 1.320 ;
        RECT  0.645 0.295 0.755 0.590 ;
        RECT  0.185 0.500 0.645 0.590 ;
        RECT  0.075 0.305 0.185 0.590 ;
    END
END OR3XD1

MACRO OR4D0
    CLASS CORE ;
    FOREIGN OR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.275 1.550 1.490 ;
        RECT  1.420 0.275 1.450 0.485 ;
        RECT  1.420 1.260 1.450 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.940 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.150 1.090 ;
        RECT  0.990 0.710 1.045 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.165 1.600 0.165 ;
        RECT  1.190 -0.165 1.300 0.410 ;
        RECT  0.680 -0.165 1.190 0.165 ;
        RECT  1.095 0.305 1.190 0.410 ;
        RECT  0.680 0.305 0.760 0.410 ;
        RECT  0.570 -0.165 0.680 0.410 ;
        RECT  0.200 -0.165 0.570 0.165 ;
        RECT  0.090 -0.165 0.200 0.475 ;
        RECT  0.000 -0.165 0.090 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.295 1.635 1.600 1.965 ;
        RECT  1.185 1.390 1.295 1.965 ;
        RECT  1.085 1.390 1.185 1.495 ;
        RECT  0.000 1.635 1.185 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.750 1.350 0.920 ;
        RECT  1.240 0.500 1.330 1.300 ;
        RECT  0.980 0.500 1.240 0.600 ;
        RECT  0.200 1.200 1.240 1.300 ;
        RECT  0.870 0.275 0.980 0.600 ;
        RECT  0.460 0.500 0.870 0.600 ;
        RECT  0.350 0.275 0.460 0.600 ;
        RECT  0.090 1.200 0.200 1.490 ;
    END
END OR4D0

MACRO OR4D1
    CLASS CORE ;
    FOREIGN OR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.310 1.550 1.490 ;
        RECT  1.420 0.310 1.450 0.600 ;
        RECT  1.420 1.060 1.450 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.940 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.150 1.090 ;
        RECT  0.990 0.710 1.045 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.165 1.600 0.165 ;
        RECT  1.190 -0.165 1.300 0.410 ;
        RECT  0.680 -0.165 1.190 0.165 ;
        RECT  1.095 0.305 1.190 0.410 ;
        RECT  0.680 0.305 0.760 0.410 ;
        RECT  0.570 -0.165 0.680 0.410 ;
        RECT  0.200 -0.165 0.570 0.165 ;
        RECT  0.090 -0.165 0.200 0.475 ;
        RECT  0.000 -0.165 0.090 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.295 1.635 1.600 1.965 ;
        RECT  1.185 1.390 1.295 1.965 ;
        RECT  1.085 1.390 1.185 1.495 ;
        RECT  0.000 1.635 1.185 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.750 1.350 0.920 ;
        RECT  1.240 0.500 1.330 1.300 ;
        RECT  0.980 0.500 1.240 0.600 ;
        RECT  0.060 1.200 1.240 1.300 ;
        RECT  0.870 0.275 0.980 0.600 ;
        RECT  0.460 0.500 0.870 0.600 ;
        RECT  0.350 0.275 0.460 0.600 ;
    END
END OR4D1

MACRO OR4D2
    CLASS CORE ;
    FOREIGN OR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.305 1.550 1.495 ;
        RECT  1.315 0.305 1.450 0.410 ;
        RECT  1.335 1.395 1.450 1.495 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0429 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.710 0.555 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0433 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.785 0.920 ;
        RECT  0.650 0.710 0.750 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  0.940 0.710 1.050 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.165 1.800 0.165 ;
        RECT  0.075 -0.165 0.185 0.485 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.635 1.800 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.500 1.340 1.305 ;
        RECT  0.995 0.500 1.240 0.600 ;
        RECT  0.060 1.200 1.240 1.305 ;
        RECT  0.885 0.325 0.995 0.600 ;
        RECT  0.295 0.325 0.885 0.435 ;
    END
END OR4D2

MACRO OR4D4
    CLASS CORE ;
    FOREIGN OR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.275 3.070 0.695 ;
        RECT  3.050 1.040 3.070 1.470 ;
        RECT  2.955 0.275 3.050 1.470 ;
        RECT  2.750 0.525 2.955 1.210 ;
        RECT  2.545 0.525 2.750 0.695 ;
        RECT  2.545 1.040 2.750 1.210 ;
        RECT  2.440 0.275 2.545 0.695 ;
        RECT  2.440 1.040 2.545 1.470 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.350 0.890 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.560 1.090 ;
        RECT  0.950 1.000 1.450 1.090 ;
        RECT  0.780 0.710 0.950 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1100 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.780 1.890 0.890 ;
        RECT  1.650 0.710 1.750 1.290 ;
        RECT  0.550 1.200 1.650 1.290 ;
        RECT  0.430 0.710 0.550 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.035 0.510 2.150 1.090 ;
        RECT  0.180 0.510 2.035 0.600 ;
        RECT  0.050 0.510 0.180 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.325 -0.165 3.400 0.165 ;
        RECT  3.215 -0.165 3.325 0.685 ;
        RECT  2.755 -0.165 3.215 0.165 ;
        RECT  2.755 0.305 2.855 0.415 ;
        RECT  2.645 -0.165 2.755 0.415 ;
        RECT  0.000 -0.165 2.645 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.325 1.635 3.400 1.965 ;
        RECT  3.215 1.050 3.325 1.965 ;
        RECT  2.805 1.635 3.215 1.965 ;
        RECT  2.695 1.300 2.805 1.965 ;
        RECT  0.185 1.635 2.695 1.965 ;
        RECT  0.075 1.050 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.545 0.525 2.650 0.695 ;
        RECT  2.545 1.040 2.650 1.210 ;
        RECT  2.440 0.275 2.545 0.695 ;
        RECT  2.440 1.040 2.545 1.470 ;
        RECT  2.350 0.785 2.595 0.890 ;
        RECT  2.260 0.310 2.350 1.490 ;
        RECT  0.285 0.310 2.260 0.420 ;
        RECT  1.065 1.380 2.260 1.490 ;
    END
END OR4D4

MACRO OR4D8
    CLASS CORE ;
    FOREIGN OR4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.955 0.275 5.065 0.685 ;
        RECT  4.955 1.050 5.065 1.460 ;
        RECT  4.565 0.585 4.955 0.685 ;
        RECT  4.565 1.050 4.955 1.150 ;
        RECT  4.455 0.275 4.565 0.685 ;
        RECT  4.455 1.050 4.565 1.460 ;
        RECT  4.250 0.585 4.455 0.685 ;
        RECT  4.250 1.050 4.455 1.150 ;
        RECT  4.045 0.585 4.250 1.150 ;
        RECT  3.950 0.275 4.045 1.460 ;
        RECT  3.935 0.275 3.950 0.685 ;
        RECT  3.935 1.050 3.950 1.460 ;
        RECT  3.525 0.585 3.935 0.685 ;
        RECT  3.525 1.050 3.935 1.150 ;
        RECT  3.415 0.275 3.525 0.685 ;
        RECT  3.415 1.050 3.525 1.460 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.700 2.955 1.100 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.700 2.155 1.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.355 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1638 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.700 0.555 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.325 -0.165 5.400 0.165 ;
        RECT  5.215 -0.165 5.325 0.685 ;
        RECT  4.305 -0.165 5.215 0.165 ;
        RECT  4.195 -0.165 4.305 0.475 ;
        RECT  3.845 -0.165 4.195 0.165 ;
        RECT  3.735 -0.165 3.845 0.475 ;
        RECT  2.305 -0.165 3.735 0.165 ;
        RECT  3.635 0.365 3.735 0.475 ;
        RECT  2.115 -0.165 2.305 0.410 ;
        RECT  1.785 -0.165 2.115 0.165 ;
        RECT  1.595 -0.165 1.785 0.410 ;
        RECT  1.265 -0.165 1.595 0.165 ;
        RECT  1.075 -0.165 1.265 0.410 ;
        RECT  0.745 -0.165 1.075 0.165 ;
        RECT  0.555 -0.165 0.745 0.410 ;
        RECT  0.185 -0.165 0.555 0.165 ;
        RECT  0.075 -0.165 0.185 0.685 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.325 1.635 5.400 1.965 ;
        RECT  5.215 1.050 5.325 1.965 ;
        RECT  4.305 1.635 5.215 1.965 ;
        RECT  4.195 1.260 4.305 1.965 ;
        RECT  3.845 1.635 4.195 1.965 ;
        RECT  3.735 1.260 3.845 1.965 ;
        RECT  3.635 1.260 3.735 1.370 ;
        RECT  0.000 1.635 3.735 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.955 0.275 5.065 0.685 ;
        RECT  4.955 1.050 5.065 1.460 ;
        RECT  4.565 0.585 4.955 0.685 ;
        RECT  4.565 1.050 4.955 1.150 ;
        RECT  4.455 0.275 4.565 0.685 ;
        RECT  4.455 1.050 4.565 1.460 ;
        RECT  4.350 0.585 4.455 0.685 ;
        RECT  4.350 1.050 4.455 1.150 ;
        RECT  3.525 0.585 3.850 0.685 ;
        RECT  3.525 1.050 3.850 1.150 ;
        RECT  3.415 0.275 3.525 0.685 ;
        RECT  3.415 1.050 3.525 1.460 ;
        RECT  3.265 0.780 3.740 0.890 ;
        RECT  3.175 0.500 3.265 0.890 ;
        RECT  2.525 0.500 3.175 0.590 ;
        RECT  2.525 1.210 3.075 1.300 ;
        RECT  2.415 0.275 2.525 0.685 ;
        RECT  2.415 1.050 2.525 1.490 ;
        RECT  0.965 0.500 2.415 0.590 ;
        RECT  1.855 1.390 2.415 1.490 ;
        RECT  1.745 1.210 2.305 1.300 ;
        RECT  1.635 1.050 1.745 1.460 ;
        RECT  1.075 1.210 1.635 1.300 ;
        RECT  0.295 1.390 1.525 1.490 ;
        RECT  0.855 0.275 0.965 1.300 ;
        RECT  0.445 0.500 0.855 0.590 ;
        RECT  0.185 1.210 0.855 1.300 ;
        RECT  0.335 0.400 0.445 0.590 ;
        RECT  0.075 1.050 0.185 1.460 ;
    END
END OR4D8

MACRO OR4XD1
    CLASS CORE ;
    FOREIGN OR4XD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1540 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.310 1.550 1.490 ;
        RECT  1.420 0.310 1.450 0.600 ;
        RECT  1.420 1.060 1.450 1.490 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.175 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.710 0.550 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.810 0.940 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.150 1.090 ;
        RECT  0.990 0.710 1.045 0.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.165 1.600 0.165 ;
        RECT  1.190 -0.165 1.300 0.410 ;
        RECT  0.680 -0.165 1.190 0.165 ;
        RECT  1.095 0.305 1.190 0.410 ;
        RECT  0.680 0.305 0.760 0.410 ;
        RECT  0.570 -0.165 0.680 0.410 ;
        RECT  0.200 -0.165 0.570 0.165 ;
        RECT  0.090 -0.165 0.200 0.475 ;
        RECT  0.000 -0.165 0.090 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.295 1.635 1.600 1.965 ;
        RECT  1.185 1.390 1.295 1.965 ;
        RECT  1.085 1.390 1.185 1.495 ;
        RECT  0.000 1.635 1.185 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.750 1.350 0.920 ;
        RECT  1.240 0.500 1.330 1.300 ;
        RECT  0.980 0.500 1.240 0.600 ;
        RECT  0.060 1.200 1.240 1.300 ;
        RECT  0.870 0.275 0.980 0.600 ;
        RECT  0.460 0.500 0.870 0.600 ;
        RECT  0.350 0.275 0.460 0.600 ;
    END
END OR4XD1

MACRO SDFCND0
    CLASS CORE ;
    FOREIGN SDFCND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.485 6.150 1.490 ;
        RECT  6.020 0.485 6.050 0.675 ;
        RECT  6.010 1.280 6.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.505 5.750 1.440 ;
        RECT  5.475 0.505 5.650 0.615 ;
        RECT  5.460 1.330 5.650 1.440 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.880 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0667 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.005 0.910 5.150 1.090 ;
        RECT  4.850 0.845 5.005 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.825 -0.165 6.200 0.165 ;
        RECT  4.655 -0.165 4.825 0.355 ;
        RECT  3.520 -0.165 4.655 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.635 6.200 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.930 0.750 5.960 0.920 ;
        RECT  5.840 0.275 5.930 0.920 ;
        RECT  5.080 0.275 5.840 0.365 ;
        RECT  5.370 0.735 5.560 0.845 ;
        RECT  5.350 1.015 5.540 1.125 ;
        RECT  5.270 0.455 5.370 0.845 ;
        RECT  5.260 1.015 5.350 1.525 ;
        RECT  5.250 0.455 5.270 0.715 ;
        RECT  4.315 1.435 5.260 1.525 ;
        RECT  4.755 0.625 5.250 0.715 ;
        RECT  4.755 1.225 5.150 1.335 ;
        RECT  4.990 0.275 5.080 0.535 ;
        RECT  4.575 0.445 4.990 0.535 ;
        RECT  4.665 0.625 4.755 1.335 ;
        RECT  4.485 0.445 4.575 1.335 ;
        RECT  4.410 0.445 4.485 0.640 ;
        RECT  4.405 1.225 4.485 1.335 ;
        RECT  4.320 0.750 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  4.230 0.315 4.285 0.840 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.665 ;
        RECT  2.390 0.565 2.585 0.665 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.565 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  0.945 1.295 2.305 1.385 ;
        RECT  2.110 0.565 2.280 0.675 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.500 1.960 1.195 ;
        RECT  1.615 0.500 1.860 0.610 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.260 0.500 1.360 0.845 ;
        RECT  0.850 0.500 1.260 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.500 0.850 0.915 ;
        RECT  0.355 0.500 0.740 0.590 ;
        RECT  0.265 0.500 0.355 1.290 ;
        RECT  0.185 0.500 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCND0

MACRO SDFCND1
    CLASS CORE ;
    FOREIGN SDFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1480 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.285 6.150 1.490 ;
        RECT  6.020 0.285 6.050 0.675 ;
        RECT  6.010 1.050 6.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.505 5.750 1.410 ;
        RECT  5.475 0.505 5.650 0.615 ;
        RECT  5.460 1.300 5.650 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0670 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.005 0.910 5.150 1.090 ;
        RECT  4.850 0.845 5.005 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.875 -0.165 6.200 0.165 ;
        RECT  4.705 -0.165 4.875 0.355 ;
        RECT  3.520 -0.165 4.705 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.635 6.200 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.930 0.750 5.960 0.920 ;
        RECT  5.840 0.275 5.930 0.920 ;
        RECT  5.080 0.275 5.840 0.365 ;
        RECT  5.370 0.735 5.560 0.845 ;
        RECT  5.370 1.015 5.540 1.125 ;
        RECT  5.270 0.455 5.370 0.845 ;
        RECT  5.280 1.015 5.370 1.525 ;
        RECT  4.315 1.435 5.280 1.525 ;
        RECT  5.250 0.455 5.270 0.715 ;
        RECT  4.755 0.625 5.250 0.715 ;
        RECT  4.755 1.225 5.150 1.335 ;
        RECT  4.990 0.275 5.080 0.535 ;
        RECT  4.575 0.445 4.990 0.535 ;
        RECT  4.665 0.625 4.755 1.335 ;
        RECT  4.485 0.445 4.575 1.335 ;
        RECT  4.410 0.445 4.485 0.625 ;
        RECT  4.405 1.225 4.485 1.335 ;
        RECT  4.320 0.730 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  4.230 0.315 4.285 0.820 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.665 ;
        RECT  2.390 0.565 2.585 0.665 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.565 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.565 2.280 0.675 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCND1

MACRO SDFCND2
    CLASS CORE ;
    FOREIGN SDFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.660 0.575 6.750 1.150 ;
        RECT  6.650 0.285 6.660 1.460 ;
        RECT  6.550 0.285 6.650 0.675 ;
        RECT  6.550 1.050 6.650 1.460 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.455 6.150 1.490 ;
        RECT  6.030 0.455 6.050 0.645 ;
        RECT  6.030 1.050 6.050 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1006 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.005 0.910 5.150 1.090 ;
        RECT  4.850 0.845 5.005 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.920 -0.165 7.000 0.165 ;
        RECT  6.810 -0.165 6.920 0.485 ;
        RECT  4.825 -0.165 6.810 0.165 ;
        RECT  4.655 -0.165 4.825 0.355 ;
        RECT  3.520 -0.165 4.655 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.920 1.635 7.000 1.965 ;
        RECT  6.810 1.250 6.920 1.965 ;
        RECT  6.400 1.635 6.810 1.965 ;
        RECT  6.290 1.050 6.400 1.965 ;
        RECT  5.880 1.635 6.290 1.965 ;
        RECT  5.770 1.090 5.880 1.965 ;
        RECT  2.610 1.635 5.770 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.440 0.780 6.540 0.890 ;
        RECT  6.350 0.275 6.440 0.890 ;
        RECT  5.080 0.275 6.350 0.365 ;
        RECT  5.620 0.750 5.960 0.920 ;
        RECT  5.510 0.625 5.620 1.500 ;
        RECT  5.360 0.625 5.510 0.715 ;
        RECT  5.250 0.455 5.360 0.715 ;
        RECT  5.250 0.825 5.360 1.525 ;
        RECT  4.755 0.625 5.250 0.715 ;
        RECT  4.315 1.435 5.250 1.525 ;
        RECT  4.755 1.225 5.150 1.335 ;
        RECT  4.990 0.275 5.080 0.535 ;
        RECT  4.575 0.445 4.990 0.535 ;
        RECT  4.665 0.625 4.755 1.335 ;
        RECT  4.485 0.445 4.575 1.335 ;
        RECT  4.410 0.445 4.485 0.625 ;
        RECT  4.405 1.225 4.485 1.335 ;
        RECT  4.320 0.730 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  4.230 0.315 4.285 0.820 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.665 ;
        RECT  2.390 0.565 2.585 0.665 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.565 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.565 2.280 0.675 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCND2

MACRO SDFCND4
    CLASS CORE ;
    FOREIGN SDFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 0.325 8.150 0.635 ;
        RECT  8.050 1.100 8.150 1.410 ;
        RECT  7.750 0.325 8.050 1.410 ;
        RECT  7.435 0.325 7.750 0.635 ;
        RECT  7.435 1.100 7.750 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.500 7.105 0.690 ;
        RECT  6.850 1.100 7.105 1.410 ;
        RECT  6.550 0.500 6.850 1.410 ;
        RECT  6.435 0.500 6.550 0.690 ;
        RECT  6.435 1.100 6.550 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1042 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.005 0.910 5.150 1.090 ;
        RECT  4.850 0.825 5.005 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.825 -0.165 8.400 0.165 ;
        RECT  4.655 -0.165 4.825 0.355 ;
        RECT  3.520 -0.165 4.655 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.635 8.400 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  0.470 1.635 2.500 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.435 0.325 7.650 0.635 ;
        RECT  7.435 1.100 7.650 1.410 ;
        RECT  6.950 0.500 7.105 0.690 ;
        RECT  6.950 1.100 7.105 1.410 ;
        RECT  6.435 0.500 6.450 0.690 ;
        RECT  6.435 1.100 6.450 1.410 ;
        RECT  7.315 0.780 7.500 0.890 ;
        RECT  7.225 0.275 7.315 0.890 ;
        RECT  6.075 0.275 7.225 0.365 ;
        RECT  6.215 0.555 6.315 1.160 ;
        RECT  6.075 0.555 6.215 0.665 ;
        RECT  6.075 1.050 6.215 1.160 ;
        RECT  5.600 0.780 6.105 0.890 ;
        RECT  5.965 0.275 6.075 0.665 ;
        RECT  5.965 1.050 6.075 1.460 ;
        RECT  5.080 0.275 5.965 0.365 ;
        RECT  5.490 0.625 5.600 1.500 ;
        RECT  5.360 0.625 5.490 0.715 ;
        RECT  5.250 0.455 5.360 0.715 ;
        RECT  5.250 0.805 5.360 1.525 ;
        RECT  4.755 0.625 5.250 0.715 ;
        RECT  4.315 1.435 5.250 1.525 ;
        RECT  4.755 1.225 5.150 1.335 ;
        RECT  4.990 0.275 5.080 0.535 ;
        RECT  4.575 0.445 4.990 0.535 ;
        RECT  4.665 0.625 4.755 1.335 ;
        RECT  4.485 0.445 4.575 1.335 ;
        RECT  4.410 0.445 4.485 0.625 ;
        RECT  4.405 1.225 4.485 1.335 ;
        RECT  4.320 0.730 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  4.230 0.315 4.285 0.820 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.645 ;
        RECT  2.390 0.545 2.585 0.645 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCND4

MACRO SDFCNQD0
    CLASS CORE ;
    FOREIGN SDFCNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0519 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.485 5.750 1.290 ;
        RECT  5.615 0.485 5.650 0.660 ;
        RECT  5.615 1.020 5.650 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.005 0.710 1.050 0.920 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0705 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 4.950 1.090 ;
        RECT  4.775 0.710 4.850 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.695 -0.165 5.800 0.165 ;
        RECT  4.525 -0.165 4.695 0.430 ;
        RECT  3.520 -0.165 4.525 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.465 1.635 5.800 1.965 ;
        RECT  5.365 1.030 5.465 1.965 ;
        RECT  2.610 1.635 5.365 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.500 0.750 5.560 0.920 ;
        RECT  5.410 0.520 5.500 0.920 ;
        RECT  5.245 0.520 5.410 0.620 ;
        RECT  5.185 0.970 5.275 1.480 ;
        RECT  5.135 0.340 5.245 0.620 ;
        RECT  5.170 0.970 5.185 1.070 ;
        RECT  4.315 1.390 5.185 1.480 ;
        RECT  5.060 0.730 5.170 1.070 ;
        RECT  4.635 0.520 5.135 0.620 ;
        RECT  4.635 1.180 5.095 1.290 ;
        RECT  4.525 0.520 4.635 1.290 ;
        RECT  4.320 0.730 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.480 ;
        RECT  4.230 0.315 4.285 0.820 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  0.945 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.250 0.495 1.355 0.875 ;
        RECT  0.850 0.495 1.250 0.595 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.495 0.850 0.930 ;
        RECT  0.355 0.495 0.740 0.590 ;
        RECT  0.265 0.495 0.355 1.290 ;
        RECT  0.185 0.495 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCNQD0

MACRO SDFCNQD1
    CLASS CORE ;
    FOREIGN SDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.285 5.750 1.490 ;
        RECT  5.615 0.285 5.650 0.665 ;
        RECT  5.615 1.050 5.650 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0702 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 4.950 1.090 ;
        RECT  4.775 0.710 4.850 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.695 -0.165 5.800 0.165 ;
        RECT  4.525 -0.165 4.695 0.430 ;
        RECT  3.520 -0.165 4.525 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.465 1.635 5.800 1.965 ;
        RECT  5.365 1.050 5.465 1.965 ;
        RECT  2.610 1.635 5.365 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.500 0.750 5.560 0.920 ;
        RECT  5.410 0.520 5.500 0.920 ;
        RECT  5.245 0.520 5.410 0.620 ;
        RECT  5.185 0.970 5.275 1.480 ;
        RECT  5.135 0.340 5.245 0.620 ;
        RECT  5.170 0.970 5.185 1.070 ;
        RECT  4.315 1.390 5.185 1.480 ;
        RECT  5.060 0.730 5.170 1.070 ;
        RECT  4.635 0.520 5.135 0.620 ;
        RECT  4.635 1.180 5.095 1.290 ;
        RECT  4.525 0.520 4.635 1.290 ;
        RECT  4.320 0.730 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.480 ;
        RECT  4.230 0.315 4.285 0.820 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCNQD1

MACRO SDFCNQD2
    CLASS CORE ;
    FOREIGN SDFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.565 6.150 1.150 ;
        RECT  6.045 0.565 6.050 0.665 ;
        RECT  6.045 1.050 6.050 1.150 ;
        RECT  5.935 0.295 6.045 0.665 ;
        RECT  5.935 1.050 6.045 1.460 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 4.950 1.090 ;
        RECT  4.800 0.710 4.850 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.305 -0.165 6.400 0.165 ;
        RECT  6.195 -0.165 6.305 0.475 ;
        RECT  5.785 -0.165 6.195 0.165 ;
        RECT  5.675 -0.165 5.785 0.485 ;
        RECT  4.760 -0.165 5.675 0.165 ;
        RECT  4.590 -0.165 4.760 0.355 ;
        RECT  3.520 -0.165 4.590 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.305 1.635 6.400 1.965 ;
        RECT  6.195 1.250 6.305 1.965 ;
        RECT  5.785 1.635 6.195 1.965 ;
        RECT  5.675 1.050 5.785 1.965 ;
        RECT  2.610 1.635 5.675 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.525 0.780 5.930 0.890 ;
        RECT  5.415 0.505 5.525 1.460 ;
        RECT  4.660 0.505 5.415 0.615 ;
        RECT  5.155 0.730 5.265 1.525 ;
        RECT  4.315 1.435 5.155 1.525 ;
        RECT  4.660 1.225 5.055 1.335 ;
        RECT  4.550 0.505 4.660 1.335 ;
        RECT  4.320 0.730 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  4.230 0.315 4.285 0.820 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCNQD2

MACRO SDFCNQD4
    CLASS CORE ;
    FOREIGN SDFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.325 6.505 0.635 ;
        RECT  6.450 1.100 6.505 1.410 ;
        RECT  6.150 0.325 6.450 1.410 ;
        RECT  5.835 0.325 6.150 0.635 ;
        RECT  5.835 1.100 6.150 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1103 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.710 4.950 1.090 ;
        RECT  4.770 0.710 4.850 0.920 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 -0.165 6.800 0.165 ;
        RECT  4.570 -0.165 4.740 0.355 ;
        RECT  3.515 -0.165 4.570 0.165 ;
        RECT  3.405 -0.165 3.515 0.415 ;
        RECT  0.520 -0.165 3.405 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.635 6.800 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  0.470 1.635 2.500 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.500 0.325 6.505 0.635 ;
        RECT  6.500 1.100 6.505 1.410 ;
        RECT  5.835 0.325 6.050 0.635 ;
        RECT  5.835 1.100 6.050 1.410 ;
        RECT  5.475 0.780 5.900 0.890 ;
        RECT  5.365 0.505 5.475 1.460 ;
        RECT  4.640 0.505 5.365 0.615 ;
        RECT  5.125 0.730 5.235 1.525 ;
        RECT  4.315 1.435 5.125 1.525 ;
        RECT  4.640 1.225 5.025 1.335 ;
        RECT  4.530 0.505 4.640 1.335 ;
        RECT  4.280 0.315 4.390 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  3.695 0.315 4.280 0.415 ;
        RECT  4.145 1.225 4.225 1.335 ;
        RECT  4.055 0.505 4.145 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.025 0.505 4.055 0.705 ;
        RECT  3.895 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.895 1.320 ;
        RECT  3.785 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.785 1.225 ;
        RECT  3.605 0.315 3.695 0.595 ;
        RECT  3.585 0.685 3.695 0.940 ;
        RECT  3.230 0.505 3.605 0.595 ;
        RECT  2.870 0.685 3.585 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.670 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.855 0.455 2.870 0.785 ;
        RECT  2.760 0.455 2.855 1.155 ;
        RECT  2.565 1.045 2.760 1.155 ;
        RECT  2.580 0.275 2.670 0.655 ;
        RECT  2.390 0.545 2.580 0.655 ;
        RECT  2.380 0.275 2.490 0.445 ;
        RECT  2.305 1.295 2.405 1.525 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.380 0.405 ;
        RECT  0.945 1.435 2.305 1.525 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.325 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.215 1.860 1.325 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCNQD4

MACRO SDFCSND0
    CLASS CORE ;
    FOREIGN SDFCSND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0646 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.710 6.150 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.825 0.475 6.950 1.330 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.530 6.550 1.295 ;
        RECT  6.260 0.530 6.450 0.640 ;
        RECT  6.260 1.185 6.450 1.295 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0355 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  1.000 0.710 1.050 0.920 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 7.000 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.620 1.635 7.000 1.965 ;
        RECT  5.450 1.400 5.620 1.965 ;
        RECT  5.050 1.635 5.450 1.965 ;
        RECT  4.880 1.405 5.050 1.965 ;
        RECT  2.610 1.635 4.880 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.645 0.275 6.735 1.515 ;
        RECT  6.105 0.275 6.645 0.375 ;
        RECT  5.910 1.405 6.645 1.515 ;
        RECT  6.240 0.750 6.350 1.095 ;
        RECT  5.760 1.005 6.240 1.095 ;
        RECT  5.995 0.275 6.105 0.490 ;
        RECT  4.860 0.275 5.995 0.365 ;
        RECT  5.800 1.185 5.910 1.515 ;
        RECT  5.710 0.455 5.760 1.095 ;
        RECT  5.660 0.455 5.710 1.290 ;
        RECT  4.950 0.455 5.660 0.565 ;
        RECT  5.620 1.005 5.660 1.290 ;
        RECT  5.165 1.180 5.620 1.290 ;
        RECT  5.440 0.710 5.530 1.090 ;
        RECT  5.045 1.000 5.440 1.090 ;
        RECT  4.955 1.000 5.045 1.305 ;
        RECT  4.510 1.215 4.955 1.305 ;
        RECT  4.770 0.275 4.860 1.125 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.410 0.980 4.510 1.305 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  0.945 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.255 0.495 1.360 0.845 ;
        RECT  0.850 0.495 1.255 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.495 0.850 0.915 ;
        RECT  0.355 0.495 0.740 0.590 ;
        RECT  0.265 0.495 0.355 1.290 ;
        RECT  0.185 0.495 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSND0

MACRO SDFCSND1
    CLASS CORE ;
    FOREIGN SDFCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0646 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.710 6.150 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.825 0.285 6.950 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.510 6.550 1.295 ;
        RECT  6.240 0.510 6.450 0.620 ;
        RECT  6.260 1.185 6.450 1.295 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 7.000 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.620 1.635 7.000 1.965 ;
        RECT  5.450 1.400 5.620 1.965 ;
        RECT  5.050 1.635 5.450 1.965 ;
        RECT  4.880 1.405 5.050 1.965 ;
        RECT  2.610 1.635 4.880 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.645 0.275 6.735 1.515 ;
        RECT  6.105 0.275 6.645 0.365 ;
        RECT  5.910 1.405 6.645 1.515 ;
        RECT  6.240 0.750 6.350 1.095 ;
        RECT  5.760 1.005 6.240 1.095 ;
        RECT  5.995 0.275 6.105 0.490 ;
        RECT  4.860 0.275 5.995 0.365 ;
        RECT  5.800 1.185 5.910 1.515 ;
        RECT  5.710 0.455 5.760 1.095 ;
        RECT  5.660 0.455 5.710 1.290 ;
        RECT  4.950 0.455 5.660 0.565 ;
        RECT  5.620 1.005 5.660 1.290 ;
        RECT  5.165 1.180 5.620 1.290 ;
        RECT  5.440 0.710 5.530 1.090 ;
        RECT  5.045 1.000 5.440 1.090 ;
        RECT  4.955 1.000 5.045 1.305 ;
        RECT  4.510 1.215 4.955 1.305 ;
        RECT  4.770 0.275 4.860 1.125 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.410 0.980 4.510 1.305 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSND1

MACRO SDFCSND2
    CLASS CORE ;
    FOREIGN SDFCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0810 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.970 0.710 6.010 0.890 ;
        RECT  5.850 0.510 5.970 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.285 7.150 1.490 ;
        RECT  6.965 0.285 7.050 0.675 ;
        RECT  6.965 1.060 7.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.550 0.465 6.575 0.675 ;
        RECT  6.550 1.030 6.575 1.240 ;
        RECT  6.450 0.465 6.550 1.240 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 7.400 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.265 1.635 7.400 1.965 ;
        RECT  6.095 1.510 6.265 1.965 ;
        RECT  5.620 1.635 6.095 1.965 ;
        RECT  5.450 1.400 5.620 1.965 ;
        RECT  5.050 1.635 5.450 1.965 ;
        RECT  4.880 1.405 5.050 1.965 ;
        RECT  2.610 1.635 4.880 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.800 0.780 6.960 0.890 ;
        RECT  6.710 0.275 6.800 1.420 ;
        RECT  6.155 0.275 6.710 0.375 ;
        RECT  5.910 1.330 6.710 1.420 ;
        RECT  6.220 0.750 6.330 1.095 ;
        RECT  5.760 1.005 6.220 1.095 ;
        RECT  5.940 0.275 6.155 0.420 ;
        RECT  4.860 0.275 5.940 0.365 ;
        RECT  5.800 1.185 5.910 1.420 ;
        RECT  5.710 0.455 5.760 1.095 ;
        RECT  5.660 0.455 5.710 1.290 ;
        RECT  4.950 0.455 5.660 0.565 ;
        RECT  5.620 1.005 5.660 1.290 ;
        RECT  5.165 1.180 5.620 1.290 ;
        RECT  5.440 0.710 5.530 1.090 ;
        RECT  5.045 1.000 5.440 1.090 ;
        RECT  4.955 1.000 5.045 1.305 ;
        RECT  4.510 1.215 4.955 1.305 ;
        RECT  4.770 0.275 4.860 1.125 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.410 0.980 4.510 1.305 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSND2

MACRO SDFCSND4
    CLASS CORE ;
    FOREIGN SDFCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0811 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.710 6.550 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.450 0.315 8.550 0.645 ;
        RECT  8.450 1.090 8.550 1.420 ;
        RECT  8.150 0.315 8.450 1.420 ;
        RECT  7.835 0.315 8.150 0.645 ;
        RECT  7.835 1.090 8.150 1.420 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.505 7.505 0.675 ;
        RECT  7.250 1.070 7.505 1.240 ;
        RECT  6.950 0.505 7.250 1.240 ;
        RECT  6.835 0.505 6.950 0.675 ;
        RECT  6.835 1.070 6.950 1.240 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0895 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.710 5.550 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.040 -0.165 8.800 0.165 ;
        RECT  4.950 -0.165 5.040 0.410 ;
        RECT  3.530 -0.165 4.950 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 1.635 8.800 1.965 ;
        RECT  6.495 1.510 6.665 1.965 ;
        RECT  5.040 1.635 6.495 1.965 ;
        RECT  4.870 1.405 5.040 1.965 ;
        RECT  2.610 1.635 4.870 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  0.470 1.635 2.500 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.835 0.315 8.050 0.645 ;
        RECT  7.835 1.090 8.050 1.420 ;
        RECT  7.350 0.505 7.505 0.675 ;
        RECT  7.350 1.070 7.505 1.240 ;
        RECT  6.835 0.505 6.850 0.675 ;
        RECT  6.835 1.070 6.850 1.240 ;
        RECT  7.700 0.780 7.920 0.890 ;
        RECT  7.610 0.275 7.700 1.420 ;
        RECT  6.495 0.275 7.610 0.375 ;
        RECT  6.330 1.330 7.610 1.420 ;
        RECT  6.640 0.730 6.745 1.095 ;
        RECT  6.150 1.005 6.640 1.095 ;
        RECT  6.385 0.275 6.495 0.585 ;
        RECT  5.220 0.275 6.385 0.365 ;
        RECT  6.220 1.185 6.330 1.420 ;
        RECT  6.130 0.485 6.150 1.095 ;
        RECT  6.040 0.485 6.130 1.270 ;
        RECT  5.415 0.485 6.040 0.595 ;
        RECT  5.155 1.160 6.040 1.270 ;
        RECT  5.800 0.710 5.910 1.070 ;
        RECT  5.160 0.980 5.800 1.070 ;
        RECT  5.130 0.275 5.220 0.610 ;
        RECT  5.050 0.710 5.160 1.070 ;
        RECT  4.860 0.520 5.130 0.610 ;
        RECT  5.045 0.980 5.050 1.070 ;
        RECT  4.955 0.980 5.045 1.305 ;
        RECT  4.510 1.215 4.955 1.305 ;
        RECT  4.770 0.440 4.860 1.125 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.410 0.980 4.510 1.305 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.525 ;
        RECT  2.280 0.545 2.390 1.145 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  0.945 1.435 2.305 1.525 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.035 2.280 1.145 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.325 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.215 1.860 1.325 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSND4

MACRO SDFCSNQD0
    CLASS CORE ;
    FOREIGN SDFCSNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0646 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.720 6.035 0.890 ;
        RECT  5.845 0.510 5.950 0.890 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.480 6.550 1.125 ;
        RECT  6.410 0.480 6.450 0.670 ;
        RECT  6.360 1.015 6.450 1.125 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.880 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0624 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.245 0.510 5.355 0.890 ;
        RECT  5.135 0.690 5.245 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 6.600 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.235 1.635 6.600 1.965 ;
        RECT  6.125 1.445 6.235 1.965 ;
        RECT  5.665 1.635 6.125 1.965 ;
        RECT  5.555 1.395 5.665 1.965 ;
        RECT  5.055 1.635 5.555 1.965 ;
        RECT  4.885 1.445 5.055 1.965 ;
        RECT  2.610 1.635 4.885 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.355 1.215 6.465 1.505 ;
        RECT  5.625 1.215 6.355 1.305 ;
        RECT  6.140 0.275 6.230 1.125 ;
        RECT  5.890 0.275 6.140 0.410 ;
        RECT  5.795 1.015 6.140 1.125 ;
        RECT  4.860 0.275 5.890 0.365 ;
        RECT  5.625 0.725 5.745 0.895 ;
        RECT  5.535 0.725 5.625 1.305 ;
        RECT  5.040 1.030 5.535 1.140 ;
        RECT  5.325 1.265 5.435 1.545 ;
        RECT  4.835 1.265 5.325 1.355 ;
        RECT  5.040 0.455 5.060 0.630 ;
        RECT  4.950 0.455 5.040 1.140 ;
        RECT  4.770 0.275 4.860 1.125 ;
        RECT  4.745 1.215 4.835 1.355 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.510 1.215 4.745 1.305 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.410 0.980 4.510 1.305 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  0.945 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.260 0.500 1.360 0.845 ;
        RECT  0.850 0.500 1.260 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.500 0.850 0.915 ;
        RECT  0.355 0.500 0.740 0.590 ;
        RECT  0.265 0.500 0.355 1.290 ;
        RECT  0.185 0.500 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSNQD0

MACRO SDFCSNQD1
    CLASS CORE ;
    FOREIGN SDFCSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0622 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0581 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.710 6.150 0.890 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.510 6.550 1.295 ;
        RECT  6.240 0.510 6.450 0.620 ;
        RECT  6.260 1.185 6.450 1.295 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0535 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 6.800 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.620 1.635 6.800 1.965 ;
        RECT  5.450 1.400 5.620 1.965 ;
        RECT  5.050 1.635 5.450 1.965 ;
        RECT  4.880 1.405 5.050 1.965 ;
        RECT  2.610 1.635 4.880 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.645 0.275 6.735 1.515 ;
        RECT  6.105 0.275 6.645 0.365 ;
        RECT  5.910 1.405 6.645 1.515 ;
        RECT  6.240 0.750 6.350 1.085 ;
        RECT  5.760 0.995 6.240 1.085 ;
        RECT  5.995 0.275 6.105 0.490 ;
        RECT  4.860 0.275 5.995 0.365 ;
        RECT  5.800 1.175 5.910 1.515 ;
        RECT  5.710 0.455 5.760 1.085 ;
        RECT  5.660 0.455 5.710 1.290 ;
        RECT  4.950 0.455 5.660 0.565 ;
        RECT  5.620 0.995 5.660 1.290 ;
        RECT  5.165 1.180 5.620 1.290 ;
        RECT  5.440 0.710 5.530 1.090 ;
        RECT  5.045 1.000 5.440 1.090 ;
        RECT  4.955 1.000 5.045 1.305 ;
        RECT  4.520 1.215 4.955 1.305 ;
        RECT  4.770 0.275 4.860 1.125 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.410 0.980 4.520 1.305 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.495 ;
        RECT  2.280 0.545 2.390 1.135 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.025 2.280 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.955 ;
        RECT  0.740 0.490 0.750 0.955 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSNQD1

MACRO SDFCSNQD2
    CLASS CORE ;
    FOREIGN SDFCSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0622 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.440 0.710 6.560 1.090 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.575 7.150 1.150 ;
        RECT  7.025 0.575 7.050 0.675 ;
        RECT  7.025 1.050 7.050 1.150 ;
        RECT  6.915 0.285 7.025 0.675 ;
        RECT  6.915 1.050 7.025 1.460 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0535 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0895 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.710 5.550 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.285 -0.165 7.400 0.165 ;
        RECT  7.175 -0.165 7.285 0.485 ;
        RECT  6.765 -0.165 7.175 0.165 ;
        RECT  6.655 -0.165 6.765 0.485 ;
        RECT  4.990 -0.165 6.655 0.165 ;
        RECT  4.880 -0.165 4.990 0.410 ;
        RECT  3.530 -0.165 4.880 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.285 1.635 7.400 1.965 ;
        RECT  7.175 1.260 7.285 1.965 ;
        RECT  6.665 1.635 7.175 1.965 ;
        RECT  6.495 1.510 6.665 1.965 ;
        RECT  6.120 1.635 6.495 1.965 ;
        RECT  5.950 1.445 6.120 1.965 ;
        RECT  5.040 1.635 5.950 1.965 ;
        RECT  4.870 1.405 5.040 1.965 ;
        RECT  2.610 1.635 4.870 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  0.470 1.635 2.500 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.710 0.730 6.820 1.355 ;
        RECT  6.130 1.265 6.710 1.355 ;
        RECT  6.330 0.305 6.535 0.415 ;
        RECT  6.220 0.275 6.330 1.175 ;
        RECT  5.220 0.275 6.220 0.365 ;
        RECT  6.030 0.485 6.130 1.355 ;
        RECT  5.375 0.485 6.030 0.595 ;
        RECT  5.155 1.160 6.030 1.270 ;
        RECT  5.800 0.710 5.910 1.070 ;
        RECT  5.160 0.980 5.800 1.070 ;
        RECT  5.130 0.275 5.220 0.610 ;
        RECT  5.050 0.710 5.160 1.070 ;
        RECT  4.860 0.520 5.130 0.610 ;
        RECT  5.045 0.980 5.050 1.070 ;
        RECT  4.955 0.980 5.045 1.305 ;
        RECT  4.520 1.215 4.955 1.305 ;
        RECT  4.770 0.520 4.860 1.125 ;
        RECT  4.710 0.520 4.770 0.615 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.600 0.440 4.710 0.615 ;
        RECT  4.575 0.730 4.680 0.905 ;
        RECT  4.510 0.730 4.575 0.820 ;
        RECT  4.410 0.980 4.520 1.305 ;
        RECT  4.420 0.315 4.510 0.820 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.525 ;
        RECT  2.280 0.545 2.390 1.145 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  0.945 1.435 2.305 1.525 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.035 2.280 1.145 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.210 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.100 1.860 1.210 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.955 ;
        RECT  0.740 0.490 0.750 0.955 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSNQD2

MACRO SDFCSNQD4
    CLASS CORE ;
    FOREIGN SDFCSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0622 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.710 6.550 0.890 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.505 7.505 0.675 ;
        RECT  7.250 1.070 7.505 1.240 ;
        RECT  6.950 0.505 7.250 1.240 ;
        RECT  6.835 0.505 6.950 0.675 ;
        RECT  6.835 1.070 6.950 1.240 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0535 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0888 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.710 5.550 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.165 7.800 0.165 ;
        RECT  4.880 -0.165 4.990 0.410 ;
        RECT  3.530 -0.165 4.880 0.165 ;
        RECT  3.410 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 1.635 7.800 1.965 ;
        RECT  6.495 1.510 6.665 1.965 ;
        RECT  5.040 1.635 6.495 1.965 ;
        RECT  4.870 1.405 5.040 1.965 ;
        RECT  2.610 1.635 4.870 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  0.470 1.635 2.500 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.350 0.505 7.505 0.675 ;
        RECT  7.350 1.070 7.505 1.240 ;
        RECT  6.835 0.505 6.850 0.675 ;
        RECT  6.835 1.070 6.850 1.240 ;
        RECT  7.610 0.275 7.700 1.420 ;
        RECT  6.495 0.275 7.610 0.375 ;
        RECT  6.330 1.330 7.610 1.420 ;
        RECT  6.640 0.730 6.745 1.085 ;
        RECT  6.150 0.995 6.640 1.085 ;
        RECT  6.385 0.275 6.495 0.485 ;
        RECT  5.220 0.275 6.385 0.365 ;
        RECT  6.220 1.175 6.330 1.420 ;
        RECT  6.130 0.485 6.150 1.085 ;
        RECT  6.040 0.485 6.130 1.270 ;
        RECT  5.425 0.485 6.040 0.595 ;
        RECT  5.155 1.160 6.040 1.270 ;
        RECT  5.800 0.710 5.910 1.070 ;
        RECT  5.160 0.980 5.800 1.070 ;
        RECT  5.130 0.275 5.220 0.610 ;
        RECT  5.050 0.710 5.160 1.070 ;
        RECT  4.860 0.520 5.130 0.610 ;
        RECT  5.045 0.980 5.050 1.070 ;
        RECT  4.955 0.980 5.045 1.305 ;
        RECT  4.520 1.215 4.955 1.305 ;
        RECT  4.770 0.520 4.860 1.125 ;
        RECT  4.710 0.520 4.770 0.615 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.600 0.440 4.710 0.615 ;
        RECT  4.575 0.730 4.680 0.905 ;
        RECT  4.510 0.730 4.575 0.820 ;
        RECT  4.410 0.980 4.520 1.305 ;
        RECT  4.420 0.315 4.510 0.820 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.890 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.485 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.875 0.685 3.605 0.785 ;
        RECT  3.385 0.910 3.485 1.295 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.675 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.585 0.275 2.675 0.655 ;
        RECT  2.390 0.545 2.585 0.655 ;
        RECT  2.385 0.275 2.495 0.445 ;
        RECT  2.305 1.295 2.405 1.525 ;
        RECT  2.280 0.545 2.390 1.145 ;
        RECT  0.865 0.305 2.385 0.405 ;
        RECT  0.945 1.435 2.305 1.525 ;
        RECT  2.110 0.545 2.280 0.655 ;
        RECT  2.065 1.035 2.280 1.145 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.325 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.215 1.860 1.325 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.955 ;
        RECT  0.740 0.490 0.750 0.955 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFCSNQD4

MACRO SDFD0
    CLASS CORE ;
    FOREIGN SDFD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0581 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.485 5.350 1.290 ;
        RECT  5.215 0.485 5.250 0.665 ;
        RECT  5.215 1.035 5.250 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.455 4.575 0.645 ;
        RECT  4.550 1.045 4.565 1.290 ;
        RECT  4.450 0.455 4.550 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.880 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.400 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 1.635 5.400 1.965 ;
        RECT  5.000 1.455 5.110 1.965 ;
        RECT  3.120 1.635 5.000 1.965 ;
        RECT  3.010 1.385 3.120 1.965 ;
        RECT  1.760 1.635 3.010 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.750 5.160 0.920 ;
        RECT  4.985 0.275 5.075 0.920 ;
        RECT  4.340 0.275 4.985 0.365 ;
        RECT  4.710 0.455 4.825 1.245 ;
        RECT  3.685 1.395 4.745 1.505 ;
        RECT  4.650 0.750 4.710 0.920 ;
        RECT  4.250 0.275 4.340 1.295 ;
        RECT  3.960 0.425 4.250 0.595 ;
        RECT  3.900 1.185 4.250 1.295 ;
        RECT  3.865 0.905 3.975 1.015 ;
        RECT  3.775 0.275 3.865 1.015 ;
        RECT  3.565 0.275 3.775 0.365 ;
        RECT  3.595 0.465 3.685 1.505 ;
        RECT  3.515 0.465 3.595 0.575 ;
        RECT  3.555 1.085 3.595 1.505 ;
        RECT  3.395 0.255 3.565 0.365 ;
        RECT  3.335 0.455 3.425 1.295 ;
        RECT  2.835 0.275 3.395 0.365 ;
        RECT  3.290 0.455 3.335 0.645 ;
        RECT  3.295 1.085 3.335 1.295 ;
        RECT  3.020 1.085 3.295 1.185 ;
        RECT  3.200 0.735 3.245 0.905 ;
        RECT  3.110 0.475 3.200 0.905 ;
        RECT  2.785 0.475 3.110 0.565 ;
        RECT  2.915 0.710 3.020 1.185 ;
        RECT  2.665 0.255 2.835 0.365 ;
        RECT  2.695 0.475 2.785 1.185 ;
        RECT  2.545 0.475 2.695 0.575 ;
        RECT  2.550 1.075 2.695 1.185 ;
        RECT  2.370 0.725 2.515 0.845 ;
        RECT  2.260 1.235 2.465 1.385 ;
        RECT  2.235 0.255 2.405 0.405 ;
        RECT  2.275 0.565 2.370 1.135 ;
        RECT  2.100 0.565 2.275 0.675 ;
        RECT  2.050 1.025 2.275 1.135 ;
        RECT  0.945 1.295 2.260 1.385 ;
        RECT  0.865 0.305 2.235 0.405 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.605 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.260 0.500 1.360 0.845 ;
        RECT  0.850 0.500 1.260 0.590 ;
        RECT  0.835 1.135 0.945 1.385 ;
        RECT  0.740 0.500 0.850 0.915 ;
        RECT  0.355 0.500 0.740 0.590 ;
        RECT  0.265 0.500 0.355 1.290 ;
        RECT  0.185 0.500 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFD0

MACRO SDFD1
    CLASS CORE ;
    FOREIGN SDFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.285 5.350 1.490 ;
        RECT  5.215 0.285 5.250 0.665 ;
        RECT  5.215 1.050 5.250 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.455 4.575 0.645 ;
        RECT  4.550 1.090 4.565 1.290 ;
        RECT  4.450 0.455 4.550 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.400 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.635 5.400 1.965 ;
        RECT  3.050 1.385 3.160 1.965 ;
        RECT  0.470 1.635 3.050 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.750 5.160 0.920 ;
        RECT  4.985 0.275 5.075 0.920 ;
        RECT  4.340 0.275 4.985 0.365 ;
        RECT  4.710 0.455 4.825 1.290 ;
        RECT  3.705 1.415 4.745 1.525 ;
        RECT  4.650 0.750 4.710 0.920 ;
        RECT  4.250 0.275 4.340 1.325 ;
        RECT  3.960 0.450 4.250 0.620 ;
        RECT  3.900 1.215 4.250 1.325 ;
        RECT  3.870 0.955 4.015 1.065 ;
        RECT  3.780 0.275 3.870 1.065 ;
        RECT  3.605 0.275 3.780 0.365 ;
        RECT  3.690 1.285 3.705 1.525 ;
        RECT  3.580 0.455 3.690 1.525 ;
        RECT  3.435 0.255 3.605 0.365 ;
        RECT  3.375 0.455 3.465 1.295 ;
        RECT  2.875 0.275 3.435 0.365 ;
        RECT  3.330 0.455 3.375 0.645 ;
        RECT  3.335 1.085 3.375 1.295 ;
        RECT  3.060 1.085 3.335 1.185 ;
        RECT  3.240 0.735 3.285 0.905 ;
        RECT  3.150 0.475 3.240 0.905 ;
        RECT  2.825 0.475 3.150 0.565 ;
        RECT  2.955 0.710 3.060 1.185 ;
        RECT  2.705 0.255 2.875 0.365 ;
        RECT  2.735 0.475 2.825 1.185 ;
        RECT  2.585 0.475 2.735 0.575 ;
        RECT  2.590 1.075 2.735 1.185 ;
        RECT  2.410 0.745 2.555 0.865 ;
        RECT  2.320 1.235 2.505 1.525 ;
        RECT  2.275 0.255 2.445 0.405 ;
        RECT  2.315 0.565 2.410 1.135 ;
        RECT  0.945 1.435 2.320 1.525 ;
        RECT  2.110 0.565 2.315 0.675 ;
        RECT  2.050 1.025 2.315 1.135 ;
        RECT  0.865 0.305 2.275 0.405 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFD1

MACRO SDFD2
    CLASS CORE ;
    FOREIGN SDFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.565 5.750 1.150 ;
        RECT  5.645 0.565 5.650 0.665 ;
        RECT  5.645 1.050 5.650 1.150 ;
        RECT  5.535 0.285 5.645 0.665 ;
        RECT  5.535 1.050 5.645 1.460 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.350 1.110 4.585 1.290 ;
        RECT  4.350 0.510 4.575 0.690 ;
        RECT  4.250 0.510 4.350 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.905 -0.165 6.000 0.165 ;
        RECT  5.795 -0.165 5.905 0.475 ;
        RECT  0.520 -0.165 5.795 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.905 1.635 6.000 1.965 ;
        RECT  5.795 1.250 5.905 1.965 ;
        RECT  5.385 1.635 5.795 1.965 ;
        RECT  5.275 1.050 5.385 1.965 ;
        RECT  3.130 1.635 5.275 1.965 ;
        RECT  3.020 1.385 3.130 1.965 ;
        RECT  0.470 1.635 3.020 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.365 0.750 5.480 0.920 ;
        RECT  5.275 0.275 5.365 0.920 ;
        RECT  4.155 0.275 5.275 0.365 ;
        RECT  5.065 0.505 5.155 1.460 ;
        RECT  4.755 0.505 5.065 0.615 ;
        RECT  5.025 1.050 5.065 1.460 ;
        RECT  4.845 0.750 4.935 1.505 ;
        RECT  3.695 1.395 4.845 1.505 ;
        RECT  4.665 0.505 4.755 0.890 ;
        RECT  4.460 0.780 4.665 0.890 ;
        RECT  4.065 0.275 4.155 1.295 ;
        RECT  3.970 0.425 4.065 0.595 ;
        RECT  3.910 1.185 4.065 1.295 ;
        RECT  3.875 0.905 3.975 1.015 ;
        RECT  3.785 0.275 3.875 1.015 ;
        RECT  3.575 0.275 3.785 0.365 ;
        RECT  3.605 0.465 3.695 1.505 ;
        RECT  3.525 0.465 3.605 0.575 ;
        RECT  3.565 1.085 3.605 1.505 ;
        RECT  3.405 0.255 3.575 0.365 ;
        RECT  3.345 0.455 3.435 1.295 ;
        RECT  2.845 0.275 3.405 0.365 ;
        RECT  3.300 0.455 3.345 0.645 ;
        RECT  3.305 1.085 3.345 1.295 ;
        RECT  3.030 1.085 3.305 1.185 ;
        RECT  3.210 0.735 3.255 0.905 ;
        RECT  3.120 0.475 3.210 0.905 ;
        RECT  2.795 0.475 3.120 0.565 ;
        RECT  2.925 0.710 3.030 1.185 ;
        RECT  2.675 0.255 2.845 0.365 ;
        RECT  2.705 0.475 2.795 1.185 ;
        RECT  2.555 0.475 2.705 0.575 ;
        RECT  2.560 1.075 2.705 1.185 ;
        RECT  2.380 0.735 2.525 0.845 ;
        RECT  2.280 1.235 2.475 1.525 ;
        RECT  2.245 0.255 2.415 0.405 ;
        RECT  2.285 0.565 2.380 1.135 ;
        RECT  2.110 0.565 2.285 0.675 ;
        RECT  2.050 1.025 2.285 1.135 ;
        RECT  0.945 1.435 2.280 1.525 ;
        RECT  0.865 0.305 2.245 0.405 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFD2

MACRO SDFD4
    CLASS CORE ;
    FOREIGN SDFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.325 7.150 0.635 ;
        RECT  7.050 1.100 7.150 1.405 ;
        RECT  6.750 0.325 7.050 1.405 ;
        RECT  6.435 0.325 6.750 0.635 ;
        RECT  6.435 1.100 6.750 1.405 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 1.100 6.150 1.410 ;
        RECT  6.050 0.520 6.105 0.690 ;
        RECT  5.750 0.520 6.050 1.410 ;
        RECT  5.435 0.520 5.750 0.690 ;
        RECT  5.435 1.100 5.750 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 7.400 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.190 1.635 7.400 1.965 ;
        RECT  3.080 1.385 3.190 1.965 ;
        RECT  0.470 1.635 3.080 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.435 0.325 6.650 0.635 ;
        RECT  6.435 1.100 6.650 1.405 ;
        RECT  5.435 0.520 5.650 0.690 ;
        RECT  5.435 1.100 5.650 1.410 ;
        RECT  6.315 0.780 6.500 0.890 ;
        RECT  6.215 0.315 6.315 0.890 ;
        RECT  4.200 0.315 6.215 0.405 ;
        RECT  5.135 0.780 5.500 0.890 ;
        RECT  5.045 0.515 5.135 1.410 ;
        RECT  4.580 0.515 5.045 0.625 ;
        RECT  4.915 1.300 5.045 1.410 ;
        RECT  4.845 0.750 4.955 1.190 ;
        RECT  4.805 1.080 4.845 1.190 ;
        RECT  4.695 1.080 4.805 1.525 ;
        RECT  3.735 1.420 4.695 1.525 ;
        RECT  4.200 1.220 4.605 1.330 ;
        RECT  4.470 0.515 4.580 0.930 ;
        RECT  4.100 0.315 4.200 1.330 ;
        RECT  3.985 0.475 4.100 0.645 ;
        RECT  3.895 1.220 4.100 1.330 ;
        RECT  3.895 0.755 3.995 1.095 ;
        RECT  3.885 0.275 3.895 1.095 ;
        RECT  3.805 0.275 3.885 0.845 ;
        RECT  3.635 0.275 3.805 0.365 ;
        RECT  3.715 1.085 3.735 1.525 ;
        RECT  3.615 0.475 3.715 1.525 ;
        RECT  3.465 0.255 3.635 0.365 ;
        RECT  3.405 0.455 3.495 1.295 ;
        RECT  2.910 0.275 3.465 0.365 ;
        RECT  3.360 0.455 3.405 0.645 ;
        RECT  3.365 1.085 3.405 1.295 ;
        RECT  3.090 1.085 3.365 1.185 ;
        RECT  3.270 0.735 3.315 0.905 ;
        RECT  3.180 0.475 3.270 0.905 ;
        RECT  2.855 0.475 3.180 0.565 ;
        RECT  2.985 0.710 3.090 1.185 ;
        RECT  2.740 0.255 2.910 0.365 ;
        RECT  2.765 0.475 2.855 1.185 ;
        RECT  2.620 0.475 2.765 0.575 ;
        RECT  2.620 1.075 2.765 1.185 ;
        RECT  2.440 0.765 2.585 0.875 ;
        RECT  2.340 1.240 2.535 1.385 ;
        RECT  2.310 0.255 2.480 0.405 ;
        RECT  2.345 0.545 2.440 1.135 ;
        RECT  2.110 0.545 2.345 0.655 ;
        RECT  2.095 1.025 2.345 1.135 ;
        RECT  1.460 1.295 2.340 1.385 ;
        RECT  0.865 0.305 2.310 0.405 ;
        RECT  1.975 0.800 2.130 0.910 ;
        RECT  1.875 0.510 1.975 1.195 ;
        RECT  1.615 0.510 1.875 0.620 ;
        RECT  1.555 1.085 1.875 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFD4

MACRO SDFKCND0
    CLASS CORE ;
    FOREIGN SDFKCND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.730 1.325 0.920 ;
        RECT  1.155 0.730 1.215 0.825 ;
        RECT  1.045 0.310 1.155 0.825 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0436 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.510 1.775 0.945 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0780 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.455 5.950 1.290 ;
        RECT  5.820 0.455 5.850 0.675 ;
        RECT  5.820 1.055 5.850 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.440 0.505 5.550 1.200 ;
        RECT  5.320 0.505 5.440 0.675 ;
        RECT  5.320 0.995 5.440 1.200 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0275 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.680 0.175 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.185 0.750 2.360 0.920 ;
        RECT  2.095 0.750 2.185 1.290 ;
        RECT  2.045 0.880 2.095 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.555 1.120 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.710 -0.165 6.000 0.165 ;
        RECT  3.710 0.465 3.930 0.585 ;
        RECT  3.600 -0.165 3.710 0.585 ;
        RECT  1.355 -0.165 3.600 0.165 ;
        RECT  1.245 -0.165 1.355 0.630 ;
        RECT  0.175 -0.165 1.245 0.165 ;
        RECT  0.065 -0.165 0.175 0.580 ;
        RECT  0.000 -0.165 0.065 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.620 1.635 6.000 1.965 ;
        RECT  3.620 1.120 3.985 1.230 ;
        RECT  3.520 1.120 3.620 1.965 ;
        RECT  1.485 1.635 3.520 1.965 ;
        RECT  1.305 1.415 1.485 1.965 ;
        RECT  0.000 1.635 1.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.730 0.775 5.755 0.945 ;
        RECT  5.640 0.775 5.730 1.495 ;
        RECT  5.230 1.375 5.640 1.495 ;
        RECT  5.160 0.600 5.230 1.495 ;
        RECT  5.140 0.300 5.160 1.495 ;
        RECT  5.050 0.300 5.140 0.710 ;
        RECT  5.045 1.380 5.140 1.495 ;
        RECT  4.670 0.600 5.050 0.710 ;
        RECT  4.880 0.830 5.050 1.000 ;
        RECT  4.790 0.830 4.880 1.495 ;
        RECT  4.580 0.830 4.790 0.920 ;
        RECT  4.300 1.380 4.790 1.495 ;
        RECT  4.390 1.100 4.650 1.230 ;
        RECT  4.480 0.295 4.580 0.920 ;
        RECT  4.310 0.295 4.480 0.425 ;
        RECT  4.280 0.550 4.390 1.230 ;
        RECT  4.090 0.300 4.190 1.515 ;
        RECT  4.070 0.300 4.090 0.565 ;
        RECT  3.715 1.345 4.090 1.515 ;
        RECT  3.890 0.675 4.000 0.910 ;
        RECT  3.430 0.675 3.890 0.765 ;
        RECT  3.380 0.675 3.430 1.280 ;
        RECT  3.315 0.275 3.380 1.280 ;
        RECT  3.270 0.275 3.315 0.765 ;
        RECT  3.065 0.275 3.165 1.495 ;
        RECT  2.200 0.275 3.065 0.405 ;
        RECT  2.010 1.395 3.065 1.495 ;
        RECT  2.870 0.510 2.975 1.170 ;
        RECT  2.695 0.510 2.870 0.640 ;
        RECT  2.725 1.060 2.870 1.170 ;
        RECT  2.575 0.750 2.740 0.920 ;
        RECT  2.475 0.545 2.575 1.200 ;
        RECT  2.215 0.545 2.475 0.655 ;
        RECT  2.275 1.030 2.475 1.200 ;
        RECT  2.010 0.265 2.200 0.405 ;
        RECT  1.955 0.595 2.005 0.790 ;
        RECT  1.865 0.595 1.955 1.305 ;
        RECT  0.955 1.215 1.865 1.305 ;
        RECT  1.555 1.035 1.720 1.125 ;
        RECT  1.555 0.295 1.675 0.420 ;
        RECT  1.445 0.295 1.555 1.125 ;
        RECT  1.075 1.010 1.445 1.125 ;
        RECT  0.945 0.915 1.075 1.125 ;
        RECT  0.855 1.215 0.955 1.485 ;
        RECT  0.855 0.455 0.910 0.635 ;
        RECT  0.835 0.455 0.855 1.485 ;
        RECT  0.765 0.455 0.835 1.305 ;
        RECT  0.355 0.460 0.675 0.570 ;
        RECT  0.355 1.295 0.675 1.465 ;
        RECT  0.265 0.460 0.355 1.465 ;
        RECT  0.065 1.295 0.265 1.465 ;
    END
END SDFKCND0

MACRO SDFKCND1
    CLASS CORE ;
    FOREIGN SDFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.730 1.325 0.920 ;
        RECT  1.155 0.730 1.215 0.825 ;
        RECT  1.045 0.310 1.155 0.825 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.510 1.775 0.945 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.845 0.285 5.950 1.495 ;
        RECT  5.820 0.285 5.845 0.675 ;
        RECT  5.820 1.055 5.845 1.495 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1410 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.440 0.285 5.550 1.200 ;
        RECT  5.320 0.285 5.440 0.675 ;
        RECT  5.320 0.995 5.440 1.200 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.680 0.175 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.185 0.750 2.360 0.920 ;
        RECT  2.095 0.750 2.185 1.290 ;
        RECT  2.045 0.880 2.095 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.555 1.120 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.710 -0.165 6.000 0.165 ;
        RECT  3.710 0.465 3.930 0.585 ;
        RECT  3.600 -0.165 3.710 0.585 ;
        RECT  1.355 -0.165 3.600 0.165 ;
        RECT  1.245 -0.165 1.355 0.630 ;
        RECT  0.175 -0.165 1.245 0.165 ;
        RECT  0.070 -0.165 0.175 0.550 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.620 1.635 6.000 1.965 ;
        RECT  3.620 1.120 3.985 1.230 ;
        RECT  3.520 1.120 3.620 1.965 ;
        RECT  1.485 1.635 3.520 1.965 ;
        RECT  1.305 1.415 1.485 1.965 ;
        RECT  0.000 1.635 1.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.730 0.775 5.755 0.945 ;
        RECT  5.640 0.775 5.730 1.495 ;
        RECT  5.230 1.375 5.640 1.495 ;
        RECT  5.165 0.600 5.230 1.495 ;
        RECT  5.140 0.300 5.165 1.495 ;
        RECT  5.050 0.300 5.140 0.710 ;
        RECT  5.045 1.380 5.140 1.495 ;
        RECT  4.670 0.600 5.050 0.710 ;
        RECT  4.880 0.830 5.050 1.000 ;
        RECT  4.790 0.830 4.880 1.495 ;
        RECT  4.580 0.830 4.790 0.920 ;
        RECT  4.300 1.380 4.790 1.495 ;
        RECT  4.390 1.100 4.650 1.230 ;
        RECT  4.480 0.295 4.580 0.920 ;
        RECT  4.310 0.295 4.480 0.425 ;
        RECT  4.280 0.550 4.390 1.230 ;
        RECT  4.090 0.300 4.190 1.515 ;
        RECT  4.070 0.300 4.090 0.565 ;
        RECT  3.715 1.345 4.090 1.515 ;
        RECT  3.890 0.675 4.000 0.910 ;
        RECT  3.430 0.675 3.890 0.765 ;
        RECT  3.380 0.675 3.430 1.280 ;
        RECT  3.315 0.275 3.380 1.280 ;
        RECT  3.270 0.275 3.315 0.765 ;
        RECT  3.065 0.290 3.165 1.495 ;
        RECT  2.125 0.290 3.065 0.400 ;
        RECT  2.010 1.395 3.065 1.495 ;
        RECT  2.870 0.520 2.975 1.170 ;
        RECT  2.705 0.520 2.870 0.630 ;
        RECT  2.725 1.060 2.870 1.170 ;
        RECT  2.575 0.750 2.740 0.920 ;
        RECT  2.475 0.520 2.575 1.200 ;
        RECT  2.225 0.520 2.475 0.630 ;
        RECT  2.275 1.030 2.475 1.200 ;
        RECT  2.015 0.290 2.125 0.480 ;
        RECT  1.955 0.595 2.005 0.790 ;
        RECT  1.865 0.595 1.955 1.305 ;
        RECT  0.955 1.215 1.865 1.305 ;
        RECT  1.555 1.035 1.720 1.125 ;
        RECT  1.555 0.295 1.675 0.420 ;
        RECT  1.445 0.295 1.555 1.125 ;
        RECT  1.075 1.010 1.445 1.125 ;
        RECT  0.945 0.915 1.075 1.125 ;
        RECT  0.855 1.215 0.955 1.485 ;
        RECT  0.855 0.455 0.910 0.635 ;
        RECT  0.835 0.455 0.855 1.485 ;
        RECT  0.765 0.455 0.835 1.305 ;
        RECT  0.355 1.295 0.675 1.465 ;
        RECT  0.525 0.325 0.655 0.590 ;
        RECT  0.355 0.480 0.525 0.590 ;
        RECT  0.265 0.480 0.355 1.465 ;
        RECT  0.065 1.295 0.265 1.465 ;
    END
END SDFKCND1

MACRO SDFKCND2
    CLASS CORE ;
    FOREIGN SDFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.730 1.325 0.920 ;
        RECT  1.155 0.730 1.215 0.825 ;
        RECT  1.045 0.310 1.155 0.825 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.510 1.775 0.945 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.255 0.535 6.350 1.170 ;
        RECT  6.245 0.295 6.255 1.490 ;
        RECT  6.135 0.295 6.245 0.665 ;
        RECT  6.125 1.045 6.245 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.610 0.285 5.755 1.125 ;
        RECT  5.565 0.985 5.610 1.125 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.680 0.175 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.185 0.750 2.360 0.920 ;
        RECT  2.095 0.750 2.185 1.290 ;
        RECT  2.045 0.880 2.095 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.555 1.120 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.515 -0.165 6.600 0.165 ;
        RECT  6.385 -0.165 6.515 0.445 ;
        RECT  5.995 -0.165 6.385 0.165 ;
        RECT  5.875 -0.165 5.995 0.675 ;
        RECT  5.475 -0.165 5.875 0.165 ;
        RECT  5.345 -0.165 5.475 0.685 ;
        RECT  4.940 -0.165 5.345 0.165 ;
        RECT  4.810 -0.165 4.940 0.460 ;
        RECT  3.710 -0.165 4.810 0.165 ;
        RECT  3.710 0.465 3.930 0.585 ;
        RECT  3.600 -0.165 3.710 0.585 ;
        RECT  1.355 -0.165 3.600 0.165 ;
        RECT  1.245 -0.165 1.355 0.630 ;
        RECT  0.175 -0.165 1.245 0.165 ;
        RECT  0.070 -0.165 0.175 0.550 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.515 1.635 6.600 1.965 ;
        RECT  6.385 1.330 6.515 1.965 ;
        RECT  5.780 1.635 6.385 1.965 ;
        RECT  5.780 1.395 6.035 1.505 ;
        RECT  5.620 1.395 5.780 1.965 ;
        RECT  5.310 1.395 5.620 1.505 ;
        RECT  3.620 1.635 5.620 1.965 ;
        RECT  3.620 1.120 3.985 1.230 ;
        RECT  3.520 1.120 3.620 1.965 ;
        RECT  1.485 1.635 3.520 1.965 ;
        RECT  1.305 1.415 1.485 1.965 ;
        RECT  0.000 1.635 1.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.990 0.770 6.155 0.900 ;
        RECT  5.895 0.770 5.990 1.305 ;
        RECT  5.245 1.215 5.895 1.305 ;
        RECT  5.220 0.300 5.245 1.305 ;
        RECT  5.140 0.300 5.220 1.520 ;
        RECT  5.095 0.300 5.140 0.710 ;
        RECT  5.090 1.215 5.140 1.520 ;
        RECT  4.670 0.600 5.095 0.710 ;
        RECT  4.930 0.830 5.050 1.000 ;
        RECT  4.840 0.830 4.930 1.495 ;
        RECT  4.580 0.830 4.840 0.920 ;
        RECT  4.300 1.380 4.840 1.495 ;
        RECT  4.390 1.100 4.650 1.230 ;
        RECT  4.480 0.295 4.580 0.920 ;
        RECT  4.310 0.295 4.480 0.425 ;
        RECT  4.280 0.550 4.390 1.230 ;
        RECT  4.090 0.300 4.190 1.515 ;
        RECT  4.070 0.300 4.090 0.565 ;
        RECT  3.715 1.345 4.090 1.515 ;
        RECT  3.890 0.675 4.000 0.910 ;
        RECT  3.430 0.675 3.890 0.765 ;
        RECT  3.380 0.675 3.430 1.280 ;
        RECT  3.315 0.275 3.380 1.280 ;
        RECT  3.270 0.275 3.315 0.765 ;
        RECT  3.065 0.290 3.165 1.525 ;
        RECT  2.125 0.290 3.065 0.400 ;
        RECT  2.010 1.395 3.065 1.525 ;
        RECT  2.870 0.520 2.975 1.220 ;
        RECT  2.705 0.520 2.870 0.630 ;
        RECT  2.765 1.030 2.870 1.220 ;
        RECT  2.575 0.750 2.740 0.920 ;
        RECT  2.475 0.520 2.575 1.200 ;
        RECT  2.225 0.520 2.475 0.630 ;
        RECT  2.275 1.030 2.475 1.200 ;
        RECT  2.015 0.290 2.125 0.495 ;
        RECT  1.955 0.595 2.005 0.790 ;
        RECT  1.865 0.595 1.955 1.305 ;
        RECT  0.955 1.215 1.865 1.305 ;
        RECT  1.555 1.035 1.720 1.125 ;
        RECT  1.555 0.295 1.675 0.420 ;
        RECT  1.445 0.295 1.555 1.125 ;
        RECT  1.075 1.010 1.445 1.125 ;
        RECT  0.945 0.915 1.075 1.125 ;
        RECT  0.855 1.215 0.955 1.485 ;
        RECT  0.855 0.455 0.910 0.635 ;
        RECT  0.835 0.455 0.855 1.485 ;
        RECT  0.765 0.455 0.835 1.305 ;
        RECT  0.355 1.295 0.675 1.465 ;
        RECT  0.525 0.325 0.655 0.590 ;
        RECT  0.355 0.480 0.525 0.590 ;
        RECT  0.265 0.480 0.355 1.465 ;
        RECT  0.065 1.295 0.265 1.465 ;
    END
END SDFKCND2

MACRO SDFKCND4
    CLASS CORE ;
    FOREIGN SDFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.730 1.325 0.920 ;
        RECT  1.155 0.730 1.215 0.825 ;
        RECT  1.045 0.310 1.155 0.825 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.510 1.775 0.945 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.945 0.295 8.075 0.675 ;
        RECT  7.945 1.020 8.075 1.470 ;
        RECT  7.850 0.525 7.945 0.675 ;
        RECT  7.850 1.020 7.945 1.190 ;
        RECT  7.555 0.525 7.850 1.190 ;
        RECT  7.550 0.295 7.555 1.490 ;
        RECT  7.425 0.295 7.550 0.675 ;
        RECT  7.425 1.020 7.550 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.945 7.075 1.115 ;
        RECT  6.905 0.295 7.035 0.710 ;
        RECT  6.850 0.540 6.905 0.710 ;
        RECT  6.550 0.540 6.850 1.115 ;
        RECT  6.515 0.540 6.550 0.710 ;
        RECT  6.345 0.945 6.550 1.115 ;
        RECT  6.385 0.295 6.515 0.710 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.680 0.175 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.185 0.710 2.545 0.890 ;
        RECT  2.095 0.710 2.185 1.290 ;
        RECT  2.045 0.880 2.095 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.555 1.120 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.335 -0.165 8.400 0.165 ;
        RECT  8.205 -0.165 8.335 0.695 ;
        RECT  7.835 -0.165 8.205 0.165 ;
        RECT  7.665 -0.165 7.835 0.425 ;
        RECT  7.295 -0.165 7.665 0.165 ;
        RECT  7.165 -0.165 7.295 0.675 ;
        RECT  6.775 -0.165 7.165 0.165 ;
        RECT  6.635 -0.165 6.775 0.450 ;
        RECT  5.760 -0.165 6.635 0.165 ;
        RECT  5.630 -0.165 5.760 0.450 ;
        RECT  4.485 -0.165 5.630 0.165 ;
        RECT  4.355 -0.165 4.485 0.625 ;
        RECT  3.860 -0.165 4.355 0.165 ;
        RECT  3.860 0.330 3.980 0.440 ;
        RECT  3.770 -0.165 3.860 0.440 ;
        RECT  1.925 -0.165 3.770 0.165 ;
        RECT  1.755 -0.165 1.925 0.420 ;
        RECT  1.355 -0.165 1.755 0.165 ;
        RECT  1.245 -0.165 1.355 0.630 ;
        RECT  0.175 -0.165 1.245 0.165 ;
        RECT  0.070 -0.165 0.175 0.550 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.335 1.635 8.400 1.965 ;
        RECT  8.205 1.035 8.335 1.965 ;
        RECT  7.815 1.635 8.205 1.965 ;
        RECT  7.685 1.325 7.815 1.965 ;
        RECT  6.980 1.635 7.685 1.965 ;
        RECT  6.980 1.385 7.335 1.500 ;
        RECT  6.820 1.385 6.980 1.965 ;
        RECT  6.605 1.385 6.820 1.500 ;
        RECT  5.730 1.635 6.820 1.965 ;
        RECT  5.590 1.250 5.730 1.965 ;
        RECT  4.435 1.635 5.590 1.965 ;
        RECT  4.265 1.215 4.435 1.965 ;
        RECT  3.925 1.635 4.265 1.965 ;
        RECT  3.745 1.215 3.925 1.965 ;
        RECT  1.485 1.635 3.745 1.965 ;
        RECT  1.305 1.415 1.485 1.965 ;
        RECT  0.000 1.635 1.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.950 0.295 8.075 0.675 ;
        RECT  7.950 1.020 8.075 1.470 ;
        RECT  7.425 0.295 7.450 0.675 ;
        RECT  7.425 1.020 7.450 1.490 ;
        RECT  6.950 0.945 7.075 1.115 ;
        RECT  6.950 0.295 7.035 0.710 ;
        RECT  6.385 0.295 6.450 0.710 ;
        RECT  6.345 0.945 6.450 1.115 ;
        RECT  7.285 0.800 7.450 0.910 ;
        RECT  7.195 0.800 7.285 1.295 ;
        RECT  6.030 1.205 7.195 1.295 ;
        RECT  5.935 0.255 6.030 1.480 ;
        RECT  5.895 0.255 5.935 0.710 ;
        RECT  5.890 1.250 5.935 1.480 ;
        RECT  5.495 0.600 5.895 0.710 ;
        RECT  5.725 0.855 5.835 1.085 ;
        RECT  5.500 0.855 5.725 0.945 ;
        RECT  5.410 0.855 5.500 1.495 ;
        RECT  5.400 0.855 5.410 0.955 ;
        RECT  4.675 1.380 5.410 1.495 ;
        RECT  5.310 0.275 5.400 0.955 ;
        RECT  5.200 1.090 5.320 1.270 ;
        RECT  5.125 0.275 5.310 0.415 ;
        RECT  5.090 0.560 5.200 1.270 ;
        RECT  4.745 0.275 5.125 0.365 ;
        RECT  4.935 0.455 5.000 0.895 ;
        RECT  4.875 0.455 4.935 1.270 ;
        RECT  4.805 0.805 4.875 1.270 ;
        RECT  4.220 0.805 4.805 0.895 ;
        RECT  4.615 0.275 4.745 0.640 ;
        RECT  4.545 1.060 4.675 1.495 ;
        RECT  4.145 0.455 4.220 1.110 ;
        RECT  4.130 0.455 4.145 1.285 ;
        RECT  4.115 0.455 4.130 0.625 ;
        RECT  4.035 1.020 4.130 1.285 ;
        RECT  3.990 0.740 4.040 0.910 ;
        RECT  3.790 1.020 4.035 1.110 ;
        RECT  3.900 0.540 3.990 0.910 ;
        RECT  3.420 0.540 3.900 0.630 ;
        RECT  3.680 0.740 3.790 1.110 ;
        RECT  3.310 0.330 3.420 1.365 ;
        RECT  3.120 0.265 3.210 1.525 ;
        RECT  2.995 0.265 3.120 0.375 ;
        RECT  2.010 1.395 3.120 1.525 ;
        RECT  2.940 0.485 3.030 1.295 ;
        RECT  2.165 0.275 2.995 0.375 ;
        RECT  2.820 0.485 2.940 0.655 ;
        RECT  2.760 1.160 2.940 1.295 ;
        RECT  2.730 0.735 2.755 1.070 ;
        RECT  2.635 0.475 2.730 1.070 ;
        RECT  2.255 0.475 2.635 0.585 ;
        RECT  2.430 0.980 2.635 1.070 ;
        RECT  2.300 0.980 2.430 1.250 ;
        RECT  2.040 0.275 2.165 0.475 ;
        RECT  1.955 0.595 2.005 0.790 ;
        RECT  1.865 0.595 1.955 1.305 ;
        RECT  0.955 1.215 1.865 1.305 ;
        RECT  1.555 1.035 1.720 1.125 ;
        RECT  1.555 0.295 1.665 0.420 ;
        RECT  1.445 0.295 1.555 1.125 ;
        RECT  1.075 1.010 1.445 1.125 ;
        RECT  0.945 0.915 1.075 1.125 ;
        RECT  0.855 1.215 0.955 1.485 ;
        RECT  0.855 0.455 0.910 0.635 ;
        RECT  0.765 0.455 0.855 1.485 ;
        RECT  0.355 1.295 0.675 1.465 ;
        RECT  0.525 0.325 0.655 0.590 ;
        RECT  0.355 0.480 0.525 0.590 ;
        RECT  0.265 0.480 0.355 1.465 ;
        RECT  0.065 1.295 0.265 1.465 ;
    END
END SDFKCND4

MACRO SDFKCNQD0
    CLASS CORE ;
    FOREIGN SDFKCNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.710 2.365 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0522 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.235 0.905 1.350 1.290 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0180 ;
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.285 5.550 1.490 ;
        RECT  5.415 0.285 5.450 0.665 ;
        RECT  5.415 1.040 5.450 1.490 ;
        RECT  5.140 0.575 5.415 0.665 ;
        RECT  5.040 0.575 5.140 0.940 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.550 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.710 2.750 1.090 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.160 1.100 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.265 -0.165 5.600 0.165 ;
        RECT  5.155 -0.165 5.265 0.465 ;
        RECT  1.310 -0.165 5.155 0.165 ;
        RECT  1.200 -0.165 1.310 0.615 ;
        RECT  0.755 -0.165 1.200 0.165 ;
        RECT  0.585 -0.165 0.755 0.295 ;
        RECT  0.000 -0.165 0.585 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 1.635 5.600 1.965 ;
        RECT  4.115 1.435 4.285 1.965 ;
        RECT  0.185 1.635 4.115 1.965 ;
        RECT  0.075 1.200 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.320 0.760 5.360 0.930 ;
        RECT  5.230 0.760 5.320 1.495 ;
        RECT  4.750 1.385 5.230 1.495 ;
        RECT  4.860 0.275 4.950 1.295 ;
        RECT  4.720 0.275 4.860 0.365 ;
        RECT  4.840 1.095 4.860 1.295 ;
        RECT  4.750 0.480 4.770 0.675 ;
        RECT  4.660 0.480 4.750 1.495 ;
        RECT  4.510 0.255 4.720 0.365 ;
        RECT  4.480 0.505 4.570 1.310 ;
        RECT  3.935 0.275 4.510 0.365 ;
        RECT  4.135 0.505 4.480 0.620 ;
        RECT  4.440 1.105 4.480 1.310 ;
        RECT  4.345 0.740 4.385 0.910 ;
        RECT  4.255 0.740 4.345 1.315 ;
        RECT  3.765 1.205 4.255 1.315 ;
        RECT  4.025 0.505 4.135 0.940 ;
        RECT  3.725 0.255 3.935 0.365 ;
        RECT  3.655 0.475 3.765 1.315 ;
        RECT  3.630 1.105 3.655 1.315 ;
        RECT  3.250 0.795 3.510 0.925 ;
        RECT  3.370 0.275 3.480 0.515 ;
        RECT  3.370 1.070 3.480 1.525 ;
        RECT  1.770 0.275 3.370 0.365 ;
        RECT  1.725 1.435 3.370 1.525 ;
        RECT  3.145 0.485 3.250 1.295 ;
        RECT  3.070 0.485 3.145 0.595 ;
        RECT  3.110 1.080 3.145 1.295 ;
        RECT  2.960 0.750 3.055 0.920 ;
        RECT  2.870 0.465 2.960 1.310 ;
        RECT  2.580 0.465 2.870 0.575 ;
        RECT  2.580 1.200 2.870 1.310 ;
        RECT  2.115 0.465 2.490 0.575 ;
        RECT  2.115 1.200 2.490 1.310 ;
        RECT  2.005 0.465 2.115 1.310 ;
        RECT  1.745 0.725 1.855 1.090 ;
        RECT  1.660 0.275 1.770 0.605 ;
        RECT  1.100 0.725 1.745 0.815 ;
        RECT  1.620 1.230 1.725 1.525 ;
        RECT  1.530 0.950 1.645 1.060 ;
        RECT  1.440 0.950 1.530 1.525 ;
        RECT  0.765 1.435 1.440 1.525 ;
        RECT  0.990 0.315 1.100 1.245 ;
        RECT  0.855 0.315 0.990 0.425 ;
        RECT  0.875 1.135 0.990 1.245 ;
        RECT  0.675 0.510 0.765 1.525 ;
        RECT  0.185 0.510 0.675 0.600 ;
        RECT  0.285 1.230 0.675 1.340 ;
        RECT  0.075 0.300 0.185 0.600 ;
    END
END SDFKCNQD0

MACRO SDFKCNQD1
    CLASS CORE ;
    FOREIGN SDFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.730 1.325 0.920 ;
        RECT  1.155 0.730 1.215 0.825 ;
        RECT  1.045 0.310 1.155 0.825 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.510 1.775 0.945 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.605 0.285 5.755 1.495 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.680 0.175 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.185 0.750 2.360 0.920 ;
        RECT  2.095 0.750 2.185 1.290 ;
        RECT  2.045 0.880 2.095 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.555 1.120 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.465 -0.165 5.800 0.165 ;
        RECT  5.355 -0.165 5.465 0.675 ;
        RECT  4.935 -0.165 5.355 0.165 ;
        RECT  4.825 -0.165 4.935 0.460 ;
        RECT  3.710 -0.165 4.825 0.165 ;
        RECT  3.710 0.465 3.930 0.585 ;
        RECT  3.600 -0.165 3.710 0.585 ;
        RECT  1.355 -0.165 3.600 0.165 ;
        RECT  1.245 -0.165 1.355 0.630 ;
        RECT  0.175 -0.165 1.245 0.165 ;
        RECT  0.070 -0.165 0.175 0.550 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.465 1.635 5.800 1.965 ;
        RECT  5.355 1.055 5.465 1.965 ;
        RECT  3.620 1.635 5.355 1.965 ;
        RECT  3.620 1.120 3.985 1.230 ;
        RECT  3.520 1.120 3.620 1.965 ;
        RECT  1.485 1.635 3.520 1.965 ;
        RECT  1.305 1.415 1.485 1.965 ;
        RECT  0.000 1.635 1.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.140 0.265 5.230 1.535 ;
        RECT  5.095 0.265 5.140 0.710 ;
        RECT  5.095 1.335 5.140 1.535 ;
        RECT  4.670 0.600 5.095 0.710 ;
        RECT  4.930 0.830 5.050 1.000 ;
        RECT  4.840 0.830 4.930 1.495 ;
        RECT  4.580 0.830 4.840 0.920 ;
        RECT  4.300 1.385 4.840 1.495 ;
        RECT  4.390 1.110 4.650 1.220 ;
        RECT  4.480 0.305 4.580 0.920 ;
        RECT  4.310 0.305 4.480 0.415 ;
        RECT  4.280 0.550 4.390 1.220 ;
        RECT  4.090 0.300 4.190 1.515 ;
        RECT  3.715 1.345 4.090 1.515 ;
        RECT  3.890 0.675 4.000 0.910 ;
        RECT  3.425 0.675 3.890 0.765 ;
        RECT  3.380 0.675 3.425 1.280 ;
        RECT  3.315 0.275 3.380 1.280 ;
        RECT  3.270 0.275 3.315 0.765 ;
        RECT  3.065 0.290 3.165 1.505 ;
        RECT  2.125 0.290 3.065 0.400 ;
        RECT  2.010 1.395 3.065 1.505 ;
        RECT  2.860 0.520 2.975 1.220 ;
        RECT  2.705 0.520 2.860 0.630 ;
        RECT  2.765 1.030 2.860 1.220 ;
        RECT  2.575 0.750 2.740 0.920 ;
        RECT  2.475 0.520 2.575 1.200 ;
        RECT  2.225 0.520 2.475 0.630 ;
        RECT  2.275 1.030 2.475 1.200 ;
        RECT  2.015 0.290 2.125 0.500 ;
        RECT  1.955 0.595 2.005 0.790 ;
        RECT  1.865 0.595 1.955 1.305 ;
        RECT  0.945 1.215 1.865 1.305 ;
        RECT  1.555 1.035 1.720 1.125 ;
        RECT  1.555 0.305 1.675 0.415 ;
        RECT  1.445 0.305 1.555 1.125 ;
        RECT  1.065 1.010 1.445 1.125 ;
        RECT  0.955 0.915 1.065 1.125 ;
        RECT  0.855 1.215 0.945 1.485 ;
        RECT  0.855 0.455 0.910 0.635 ;
        RECT  0.765 0.455 0.855 1.485 ;
        RECT  0.355 1.295 0.675 1.465 ;
        RECT  0.525 0.325 0.655 0.590 ;
        RECT  0.355 0.480 0.525 0.590 ;
        RECT  0.265 0.480 0.355 1.465 ;
        RECT  0.065 1.295 0.265 1.465 ;
    END
END SDFKCNQD1

MACRO SDFKCNQD2
    CLASS CORE ;
    FOREIGN SDFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.730 1.325 0.920 ;
        RECT  1.155 0.730 1.215 0.825 ;
        RECT  1.045 0.310 1.155 0.825 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.510 1.775 0.945 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.560 0.285 5.750 1.515 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.680 0.175 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.185 0.750 2.360 0.920 ;
        RECT  2.095 0.750 2.185 1.290 ;
        RECT  2.045 0.880 2.095 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.555 1.120 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.940 -0.165 6.000 0.165 ;
        RECT  4.810 -0.165 4.940 0.460 ;
        RECT  3.710 -0.165 4.810 0.165 ;
        RECT  3.710 0.465 3.930 0.585 ;
        RECT  3.600 -0.165 3.710 0.585 ;
        RECT  1.355 -0.165 3.600 0.165 ;
        RECT  1.245 -0.165 1.355 0.630 ;
        RECT  0.175 -0.165 1.245 0.165 ;
        RECT  0.070 -0.165 0.175 0.550 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.620 1.635 6.000 1.965 ;
        RECT  3.620 1.120 3.985 1.230 ;
        RECT  3.520 1.120 3.620 1.965 ;
        RECT  1.485 1.635 3.520 1.965 ;
        RECT  1.305 1.415 1.485 1.965 ;
        RECT  0.000 1.635 1.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.140 0.275 5.245 1.530 ;
        RECT  5.095 0.275 5.140 0.710 ;
        RECT  5.085 1.335 5.140 1.530 ;
        RECT  4.670 0.600 5.095 0.710 ;
        RECT  4.930 0.830 5.050 1.000 ;
        RECT  4.840 0.830 4.930 1.495 ;
        RECT  4.580 0.830 4.840 0.920 ;
        RECT  4.300 1.380 4.840 1.495 ;
        RECT  4.390 1.100 4.650 1.230 ;
        RECT  4.480 0.295 4.580 0.920 ;
        RECT  4.310 0.295 4.480 0.425 ;
        RECT  4.280 0.550 4.390 1.230 ;
        RECT  4.090 0.300 4.190 1.515 ;
        RECT  4.070 0.300 4.090 0.565 ;
        RECT  3.715 1.345 4.090 1.515 ;
        RECT  3.890 0.675 4.000 0.910 ;
        RECT  3.430 0.675 3.890 0.765 ;
        RECT  3.380 0.675 3.430 1.280 ;
        RECT  3.315 0.275 3.380 1.280 ;
        RECT  3.270 0.275 3.315 0.765 ;
        RECT  3.065 0.290 3.165 1.525 ;
        RECT  2.125 0.290 3.065 0.400 ;
        RECT  2.010 1.395 3.065 1.525 ;
        RECT  2.860 0.520 2.975 1.220 ;
        RECT  2.705 0.520 2.860 0.630 ;
        RECT  2.765 1.030 2.860 1.220 ;
        RECT  2.575 0.750 2.740 0.920 ;
        RECT  2.475 0.520 2.575 1.200 ;
        RECT  2.225 0.520 2.475 0.630 ;
        RECT  2.275 1.030 2.475 1.200 ;
        RECT  2.015 0.290 2.125 0.500 ;
        RECT  1.955 0.595 2.005 0.790 ;
        RECT  1.865 0.595 1.955 1.305 ;
        RECT  0.955 1.215 1.865 1.305 ;
        RECT  1.555 1.035 1.720 1.125 ;
        RECT  1.555 0.295 1.675 0.420 ;
        RECT  1.445 0.295 1.555 1.125 ;
        RECT  1.075 1.010 1.445 1.125 ;
        RECT  0.945 0.915 1.075 1.125 ;
        RECT  0.855 1.215 0.955 1.485 ;
        RECT  0.855 0.455 0.910 0.635 ;
        RECT  0.765 0.455 0.855 1.485 ;
        RECT  0.355 1.295 0.675 1.465 ;
        RECT  0.525 0.325 0.655 0.590 ;
        RECT  0.355 0.480 0.525 0.590 ;
        RECT  0.265 0.480 0.355 1.465 ;
        RECT  0.065 1.295 0.265 1.465 ;
    END
END SDFKCNQD2

MACRO SDFKCNQD4
    CLASS CORE ;
    FOREIGN SDFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.730 1.325 0.920 ;
        RECT  1.155 0.730 1.215 0.825 ;
        RECT  1.045 0.310 1.155 0.825 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0549 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.510 1.775 0.945 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.930 0.295 7.060 0.675 ;
        RECT  6.930 1.020 7.060 1.470 ;
        RECT  6.850 0.525 6.930 0.675 ;
        RECT  6.850 1.020 6.930 1.190 ;
        RECT  6.550 0.525 6.850 1.190 ;
        RECT  6.540 0.525 6.550 0.675 ;
        RECT  6.540 1.020 6.550 1.190 ;
        RECT  6.410 0.295 6.540 0.675 ;
        RECT  6.410 1.020 6.540 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.680 0.175 1.120 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.185 0.710 2.545 0.890 ;
        RECT  2.095 0.710 2.185 1.290 ;
        RECT  2.045 0.880 2.095 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0556 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.710 0.555 1.120 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.320 -0.165 7.400 0.165 ;
        RECT  7.190 -0.165 7.320 0.695 ;
        RECT  6.820 -0.165 7.190 0.165 ;
        RECT  6.650 -0.165 6.820 0.425 ;
        RECT  6.280 -0.165 6.650 0.165 ;
        RECT  6.150 -0.165 6.280 0.690 ;
        RECT  5.760 -0.165 6.150 0.165 ;
        RECT  5.630 -0.165 5.760 0.450 ;
        RECT  4.475 -0.165 5.630 0.165 ;
        RECT  4.365 -0.165 4.475 0.625 ;
        RECT  3.860 -0.165 4.365 0.165 ;
        RECT  3.860 0.365 3.980 0.475 ;
        RECT  3.770 -0.165 3.860 0.475 ;
        RECT  1.925 -0.165 3.770 0.165 ;
        RECT  1.755 -0.165 1.925 0.420 ;
        RECT  1.355 -0.165 1.755 0.165 ;
        RECT  1.245 -0.165 1.355 0.630 ;
        RECT  0.175 -0.165 1.245 0.165 ;
        RECT  0.070 -0.165 0.175 0.550 ;
        RECT  0.000 -0.165 0.070 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.320 1.635 7.400 1.965 ;
        RECT  7.190 1.035 7.320 1.965 ;
        RECT  6.800 1.635 7.190 1.965 ;
        RECT  6.670 1.325 6.800 1.965 ;
        RECT  6.280 1.635 6.670 1.965 ;
        RECT  6.150 1.030 6.280 1.965 ;
        RECT  5.715 1.635 6.150 1.965 ;
        RECT  5.605 1.330 5.715 1.965 ;
        RECT  4.435 1.635 5.605 1.965 ;
        RECT  4.265 1.215 4.435 1.965 ;
        RECT  3.925 1.635 4.265 1.965 ;
        RECT  3.745 1.215 3.925 1.965 ;
        RECT  1.485 1.635 3.745 1.965 ;
        RECT  1.305 1.415 1.485 1.965 ;
        RECT  0.000 1.635 1.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.950 0.295 7.060 0.675 ;
        RECT  6.950 1.020 7.060 1.470 ;
        RECT  6.410 0.295 6.450 0.675 ;
        RECT  6.410 1.020 6.450 1.490 ;
        RECT  5.935 0.255 6.030 1.525 ;
        RECT  5.895 0.255 5.935 0.710 ;
        RECT  5.890 1.335 5.935 1.525 ;
        RECT  5.495 0.600 5.895 0.710 ;
        RECT  5.725 0.855 5.835 1.085 ;
        RECT  5.500 0.855 5.725 0.945 ;
        RECT  5.410 0.855 5.500 1.495 ;
        RECT  5.400 0.855 5.410 0.955 ;
        RECT  4.665 1.385 5.410 1.495 ;
        RECT  5.310 0.275 5.400 0.955 ;
        RECT  5.205 1.090 5.320 1.270 ;
        RECT  5.125 0.275 5.310 0.415 ;
        RECT  5.095 0.560 5.205 1.270 ;
        RECT  4.735 0.275 5.125 0.365 ;
        RECT  4.925 0.455 4.995 0.895 ;
        RECT  4.885 0.455 4.925 1.270 ;
        RECT  4.815 0.805 4.885 1.270 ;
        RECT  4.220 0.805 4.815 0.895 ;
        RECT  4.625 0.275 4.735 0.640 ;
        RECT  4.555 1.060 4.665 1.495 ;
        RECT  4.145 0.455 4.220 1.110 ;
        RECT  4.130 0.455 4.145 1.285 ;
        RECT  4.105 0.455 4.130 0.625 ;
        RECT  4.035 1.020 4.130 1.285 ;
        RECT  3.990 0.740 4.040 0.910 ;
        RECT  3.790 1.020 4.035 1.110 ;
        RECT  3.900 0.575 3.990 0.910 ;
        RECT  3.420 0.575 3.900 0.665 ;
        RECT  3.680 0.775 3.790 1.110 ;
        RECT  3.310 0.330 3.420 1.365 ;
        RECT  3.120 0.265 3.210 1.525 ;
        RECT  2.995 0.265 3.120 0.375 ;
        RECT  2.010 1.395 3.120 1.525 ;
        RECT  2.940 0.485 3.030 1.275 ;
        RECT  2.155 0.275 2.995 0.375 ;
        RECT  2.820 0.485 2.940 0.655 ;
        RECT  2.760 1.165 2.940 1.275 ;
        RECT  2.730 0.735 2.755 1.070 ;
        RECT  2.635 0.475 2.730 1.070 ;
        RECT  2.255 0.475 2.635 0.585 ;
        RECT  2.420 0.980 2.635 1.070 ;
        RECT  2.310 0.980 2.420 1.250 ;
        RECT  2.045 0.275 2.155 0.475 ;
        RECT  1.955 0.595 2.005 0.790 ;
        RECT  1.865 0.595 1.955 1.305 ;
        RECT  0.945 1.215 1.865 1.305 ;
        RECT  1.555 1.035 1.720 1.125 ;
        RECT  1.555 0.305 1.665 0.415 ;
        RECT  1.445 0.305 1.555 1.125 ;
        RECT  1.065 1.010 1.445 1.125 ;
        RECT  0.955 0.915 1.065 1.125 ;
        RECT  0.855 1.215 0.945 1.485 ;
        RECT  0.855 0.455 0.905 0.635 ;
        RECT  0.835 0.455 0.855 1.485 ;
        RECT  0.765 0.455 0.835 1.305 ;
        RECT  0.355 1.295 0.675 1.465 ;
        RECT  0.535 0.325 0.645 0.590 ;
        RECT  0.355 0.480 0.535 0.590 ;
        RECT  0.265 0.480 0.355 1.465 ;
        RECT  0.065 1.295 0.265 1.465 ;
    END
END SDFKCNQD4

MACRO SDFKCSND0
    CLASS CORE ;
    FOREIGN SDFKCSND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.500 2.150 0.930 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0481 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.275 2.755 0.690 ;
        RECT  2.415 0.275 2.635 0.440 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.645 0.465 6.750 1.290 ;
        RECT  6.615 0.465 6.645 0.665 ;
        RECT  6.625 1.060 6.645 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.245 0.505 6.355 1.210 ;
        RECT  6.120 0.505 6.245 0.685 ;
        RECT  6.120 1.040 6.245 1.210 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.065 0.880 1.175 ;
        RECT  0.650 1.065 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.710 3.320 0.890 ;
        RECT  2.895 0.710 2.995 1.290 ;
        RECT  2.845 1.060 2.895 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.685 1.350 1.195 ;
        RECT  0.630 0.685 1.250 0.775 ;
        RECT  0.990 1.085 1.250 1.195 ;
        RECT  0.460 0.660 0.630 0.775 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.720 -0.165 6.800 0.165 ;
        RECT  5.610 -0.165 5.720 0.450 ;
        RECT  4.610 -0.165 5.610 0.165 ;
        RECT  4.610 0.385 4.730 0.495 ;
        RECT  4.520 -0.165 4.610 0.495 ;
        RECT  2.270 -0.165 4.520 0.165 ;
        RECT  2.160 -0.165 2.270 0.395 ;
        RECT  0.000 -0.165 2.160 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 1.635 6.800 1.965 ;
        RECT  5.575 1.250 5.685 1.965 ;
        RECT  4.675 1.635 5.575 1.965 ;
        RECT  4.495 1.215 4.675 1.965 ;
        RECT  2.685 1.635 4.495 1.965 ;
        RECT  2.555 1.440 2.685 1.965 ;
        RECT  2.300 1.635 2.555 1.965 ;
        RECT  2.130 1.415 2.300 1.965 ;
        RECT  1.260 1.635 2.130 1.965 ;
        RECT  1.090 1.495 1.260 1.965 ;
        RECT  0.500 1.635 1.090 1.965 ;
        RECT  0.330 1.495 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.535 0.775 6.555 0.945 ;
        RECT  6.445 0.775 6.535 1.410 ;
        RECT  5.995 1.320 6.445 1.410 ;
        RECT  5.955 0.265 6.055 0.365 ;
        RECT  5.970 0.600 5.995 1.410 ;
        RECT  5.955 0.600 5.970 1.545 ;
        RECT  5.905 0.265 5.955 1.545 ;
        RECT  5.865 0.265 5.905 0.710 ;
        RECT  5.860 1.320 5.905 1.545 ;
        RECT  5.465 0.600 5.865 0.710 ;
        RECT  5.695 0.855 5.805 1.085 ;
        RECT  5.470 0.855 5.695 0.945 ;
        RECT  5.380 0.855 5.470 1.495 ;
        RECT  5.370 0.855 5.380 0.955 ;
        RECT  4.995 1.385 5.380 1.495 ;
        RECT  5.280 0.305 5.370 0.955 ;
        RECT  5.170 1.090 5.290 1.270 ;
        RECT  5.090 0.305 5.280 0.415 ;
        RECT  5.060 0.560 5.170 1.270 ;
        RECT  4.895 0.465 4.970 1.110 ;
        RECT  4.880 0.465 4.895 1.285 ;
        RECT  4.865 0.465 4.880 0.635 ;
        RECT  4.785 1.020 4.880 1.285 ;
        RECT  4.740 0.740 4.790 0.910 ;
        RECT  4.540 1.020 4.785 1.110 ;
        RECT  4.650 0.595 4.740 0.910 ;
        RECT  4.170 0.595 4.650 0.685 ;
        RECT  4.430 0.795 4.540 1.110 ;
        RECT  4.060 0.330 4.170 1.365 ;
        RECT  3.870 0.265 3.960 1.525 ;
        RECT  3.745 0.265 3.870 0.375 ;
        RECT  3.050 1.435 3.870 1.525 ;
        RECT  3.680 0.485 3.780 1.275 ;
        RECT  3.035 0.275 3.745 0.375 ;
        RECT  3.595 0.485 3.680 0.655 ;
        RECT  3.535 1.165 3.680 1.275 ;
        RECT  3.505 0.735 3.530 1.070 ;
        RECT  3.410 0.510 3.505 1.070 ;
        RECT  3.055 0.510 3.410 0.620 ;
        RECT  3.195 0.980 3.410 1.070 ;
        RECT  3.085 0.980 3.195 1.250 ;
        RECT  2.835 1.415 3.050 1.525 ;
        RECT  2.845 0.265 3.035 0.375 ;
        RECT  2.700 0.780 2.805 0.950 ;
        RECT  2.610 0.780 2.700 1.320 ;
        RECT  1.760 1.230 2.610 1.320 ;
        RECT  2.370 1.030 2.510 1.140 ;
        RECT  2.370 0.545 2.490 0.655 ;
        RECT  2.260 0.545 2.370 1.140 ;
        RECT  1.910 1.035 2.260 1.140 ;
        RECT  1.800 0.885 1.910 1.140 ;
        RECT  1.710 0.480 1.835 0.595 ;
        RECT  1.710 1.230 1.760 1.475 ;
        RECT  1.620 0.480 1.710 1.475 ;
        RECT  1.440 0.390 1.530 1.395 ;
        RECT  1.415 0.390 1.440 0.595 ;
        RECT  0.945 1.305 1.440 1.395 ;
        RECT  0.830 0.495 1.415 0.595 ;
        RECT  0.695 0.295 1.295 0.405 ;
        RECT  0.560 0.865 1.140 0.975 ;
        RECT  0.840 1.305 0.945 1.495 ;
        RECT  0.585 0.295 0.695 0.510 ;
        RECT  0.440 0.865 0.560 1.195 ;
        RECT  0.350 0.865 0.440 0.965 ;
        RECT  0.260 0.500 0.350 1.385 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.045 1.275 0.260 1.385 ;
        RECT  0.075 0.300 0.185 0.590 ;
    END
END SDFKCSND0

MACRO SDFKCSND1
    CLASS CORE ;
    FOREIGN SDFKCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.500 2.150 0.930 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0539 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.275 2.755 0.690 ;
        RECT  2.415 0.275 2.635 0.440 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.645 0.295 6.750 1.490 ;
        RECT  6.615 0.295 6.645 0.665 ;
        RECT  6.625 1.060 6.645 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.245 0.505 6.355 1.210 ;
        RECT  6.120 0.505 6.245 0.685 ;
        RECT  6.120 1.040 6.245 1.210 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.065 0.880 1.175 ;
        RECT  0.650 1.065 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.710 3.320 0.890 ;
        RECT  2.895 0.710 2.995 1.290 ;
        RECT  2.845 1.060 2.895 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.685 1.350 1.215 ;
        RECT  0.630 0.685 1.250 0.775 ;
        RECT  0.990 1.105 1.250 1.215 ;
        RECT  0.460 0.660 0.630 0.775 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 -0.165 6.800 0.165 ;
        RECT  5.600 -0.165 5.730 0.450 ;
        RECT  4.610 -0.165 5.600 0.165 ;
        RECT  4.610 0.385 4.730 0.495 ;
        RECT  4.520 -0.165 4.610 0.495 ;
        RECT  2.270 -0.165 4.520 0.165 ;
        RECT  2.160 -0.165 2.270 0.395 ;
        RECT  0.000 -0.165 2.160 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 1.635 6.800 1.965 ;
        RECT  5.575 1.250 5.685 1.965 ;
        RECT  4.675 1.635 5.575 1.965 ;
        RECT  4.495 1.215 4.675 1.965 ;
        RECT  2.685 1.635 4.495 1.965 ;
        RECT  2.555 1.440 2.685 1.965 ;
        RECT  2.300 1.635 2.555 1.965 ;
        RECT  2.130 1.415 2.300 1.965 ;
        RECT  1.260 1.635 2.130 1.965 ;
        RECT  1.090 1.495 1.260 1.965 ;
        RECT  0.500 1.635 1.090 1.965 ;
        RECT  0.330 1.495 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.535 0.775 6.555 0.945 ;
        RECT  6.445 0.775 6.535 1.410 ;
        RECT  5.995 1.320 6.445 1.410 ;
        RECT  5.955 0.265 6.055 0.365 ;
        RECT  5.970 0.600 5.995 1.410 ;
        RECT  5.955 0.600 5.970 1.545 ;
        RECT  5.905 0.265 5.955 1.545 ;
        RECT  5.865 0.265 5.905 0.710 ;
        RECT  5.860 1.320 5.905 1.545 ;
        RECT  5.465 0.600 5.865 0.710 ;
        RECT  5.695 0.855 5.805 1.085 ;
        RECT  5.470 0.855 5.695 0.945 ;
        RECT  5.380 0.855 5.470 1.495 ;
        RECT  5.370 0.855 5.380 0.955 ;
        RECT  4.995 1.385 5.380 1.495 ;
        RECT  5.280 0.305 5.370 0.955 ;
        RECT  5.170 1.090 5.290 1.270 ;
        RECT  5.090 0.305 5.280 0.415 ;
        RECT  5.060 0.560 5.170 1.270 ;
        RECT  4.895 0.465 4.970 1.110 ;
        RECT  4.880 0.465 4.895 1.285 ;
        RECT  4.865 0.465 4.880 0.635 ;
        RECT  4.785 1.020 4.880 1.285 ;
        RECT  4.740 0.740 4.790 0.910 ;
        RECT  4.540 1.020 4.785 1.110 ;
        RECT  4.650 0.595 4.740 0.910 ;
        RECT  4.170 0.595 4.650 0.685 ;
        RECT  4.430 0.795 4.540 1.110 ;
        RECT  4.060 0.330 4.170 1.365 ;
        RECT  3.870 0.265 3.960 1.525 ;
        RECT  3.745 0.265 3.870 0.375 ;
        RECT  3.050 1.435 3.870 1.525 ;
        RECT  3.690 0.485 3.780 1.275 ;
        RECT  3.035 0.275 3.745 0.375 ;
        RECT  3.595 0.485 3.690 0.655 ;
        RECT  3.535 1.165 3.690 1.275 ;
        RECT  3.505 0.735 3.530 1.070 ;
        RECT  3.410 0.510 3.505 1.070 ;
        RECT  3.055 0.510 3.410 0.620 ;
        RECT  3.195 0.980 3.410 1.070 ;
        RECT  3.085 0.980 3.195 1.250 ;
        RECT  2.835 1.415 3.050 1.525 ;
        RECT  2.845 0.265 3.035 0.375 ;
        RECT  2.700 0.780 2.805 0.950 ;
        RECT  2.610 0.780 2.700 1.320 ;
        RECT  1.750 1.230 2.610 1.320 ;
        RECT  2.370 1.030 2.510 1.140 ;
        RECT  2.370 0.545 2.490 0.655 ;
        RECT  2.260 0.545 2.370 1.140 ;
        RECT  1.910 1.035 2.260 1.140 ;
        RECT  1.800 0.885 1.910 1.140 ;
        RECT  1.710 0.485 1.835 0.595 ;
        RECT  1.710 1.230 1.750 1.475 ;
        RECT  1.620 0.485 1.710 1.475 ;
        RECT  1.440 0.390 1.530 1.395 ;
        RECT  1.405 0.390 1.440 0.595 ;
        RECT  0.945 1.305 1.440 1.395 ;
        RECT  0.830 0.495 1.405 0.595 ;
        RECT  0.695 0.295 1.295 0.405 ;
        RECT  0.560 0.865 1.140 0.975 ;
        RECT  0.840 1.305 0.945 1.495 ;
        RECT  0.585 0.295 0.695 0.505 ;
        RECT  0.440 0.865 0.560 1.195 ;
        RECT  0.350 0.865 0.440 0.965 ;
        RECT  0.260 0.500 0.350 1.385 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.275 0.260 1.385 ;
        RECT  0.075 0.280 0.185 0.590 ;
        RECT  0.075 1.275 0.185 1.465 ;
    END
END SDFKCSND1

MACRO SDFKCSND2
    CLASS CORE ;
    FOREIGN SDFKCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.500 2.150 0.930 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0539 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.275 2.755 0.690 ;
        RECT  2.415 0.275 2.635 0.440 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.045 0.535 7.150 1.170 ;
        RECT  7.030 0.535 7.045 0.665 ;
        RECT  7.030 1.045 7.045 1.170 ;
        RECT  6.910 0.295 7.030 0.665 ;
        RECT  6.900 1.045 7.030 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.385 0.285 6.555 1.125 ;
        RECT  6.340 0.985 6.385 1.125 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.065 0.880 1.175 ;
        RECT  0.650 1.065 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.710 3.320 0.890 ;
        RECT  2.895 0.710 2.995 1.290 ;
        RECT  2.845 1.060 2.895 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.685 1.350 1.215 ;
        RECT  0.630 0.685 1.250 0.775 ;
        RECT  0.990 1.105 1.250 1.215 ;
        RECT  0.460 0.660 0.630 0.775 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.290 -0.165 7.400 0.165 ;
        RECT  7.160 -0.165 7.290 0.445 ;
        RECT  6.770 -0.165 7.160 0.165 ;
        RECT  6.650 -0.165 6.770 0.675 ;
        RECT  6.250 -0.165 6.650 0.165 ;
        RECT  6.120 -0.165 6.250 0.685 ;
        RECT  5.730 -0.165 6.120 0.165 ;
        RECT  5.600 -0.165 5.730 0.450 ;
        RECT  4.610 -0.165 5.600 0.165 ;
        RECT  4.610 0.385 4.730 0.495 ;
        RECT  4.520 -0.165 4.610 0.495 ;
        RECT  2.270 -0.165 4.520 0.165 ;
        RECT  2.150 -0.165 2.270 0.395 ;
        RECT  0.000 -0.165 2.150 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.285 1.635 7.400 1.965 ;
        RECT  7.170 1.330 7.285 1.965 ;
        RECT  6.580 1.635 7.170 1.965 ;
        RECT  6.580 1.395 6.810 1.505 ;
        RECT  6.420 1.395 6.580 1.965 ;
        RECT  6.085 1.395 6.420 1.505 ;
        RECT  5.700 1.635 6.420 1.965 ;
        RECT  5.560 1.250 5.700 1.965 ;
        RECT  4.675 1.635 5.560 1.965 ;
        RECT  4.495 1.215 4.675 1.965 ;
        RECT  2.685 1.635 4.495 1.965 ;
        RECT  2.555 1.440 2.685 1.965 ;
        RECT  2.300 1.635 2.555 1.965 ;
        RECT  2.130 1.415 2.300 1.965 ;
        RECT  1.260 1.635 2.130 1.965 ;
        RECT  1.090 1.495 1.260 1.965 ;
        RECT  0.500 1.635 1.090 1.965 ;
        RECT  0.330 1.495 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.765 0.770 6.935 0.920 ;
        RECT  6.670 0.770 6.765 1.305 ;
        RECT  6.015 1.215 6.670 1.305 ;
        RECT  5.995 0.255 6.015 1.305 ;
        RECT  5.905 0.255 5.995 1.480 ;
        RECT  5.865 0.255 5.905 0.710 ;
        RECT  5.860 1.250 5.905 1.480 ;
        RECT  5.465 0.600 5.865 0.710 ;
        RECT  5.695 0.855 5.805 1.085 ;
        RECT  5.470 0.855 5.695 0.945 ;
        RECT  5.380 0.855 5.470 1.495 ;
        RECT  5.370 0.855 5.380 0.955 ;
        RECT  4.995 1.380 5.380 1.495 ;
        RECT  5.280 0.305 5.370 0.955 ;
        RECT  5.170 1.090 5.290 1.270 ;
        RECT  5.090 0.305 5.280 0.415 ;
        RECT  5.060 0.560 5.170 1.270 ;
        RECT  4.895 0.465 4.970 1.110 ;
        RECT  4.880 0.465 4.895 1.285 ;
        RECT  4.865 0.465 4.880 0.635 ;
        RECT  4.785 1.020 4.880 1.285 ;
        RECT  4.740 0.740 4.790 0.910 ;
        RECT  4.540 1.020 4.785 1.110 ;
        RECT  4.650 0.595 4.740 0.910 ;
        RECT  4.170 0.595 4.650 0.685 ;
        RECT  4.430 0.795 4.540 1.110 ;
        RECT  4.060 0.330 4.170 1.365 ;
        RECT  3.870 0.265 3.960 1.525 ;
        RECT  3.745 0.265 3.870 0.375 ;
        RECT  3.050 1.435 3.870 1.525 ;
        RECT  3.690 0.485 3.780 1.295 ;
        RECT  3.035 0.275 3.745 0.375 ;
        RECT  3.595 0.485 3.690 0.655 ;
        RECT  3.535 1.160 3.690 1.295 ;
        RECT  3.505 0.735 3.530 1.070 ;
        RECT  3.410 0.510 3.505 1.070 ;
        RECT  3.055 0.510 3.410 0.620 ;
        RECT  3.195 0.980 3.410 1.070 ;
        RECT  3.085 0.980 3.195 1.250 ;
        RECT  2.835 1.415 3.050 1.525 ;
        RECT  2.845 0.265 3.035 0.375 ;
        RECT  2.700 0.780 2.805 0.950 ;
        RECT  2.610 0.780 2.700 1.320 ;
        RECT  1.760 1.230 2.610 1.320 ;
        RECT  2.370 1.030 2.510 1.140 ;
        RECT  2.370 0.530 2.490 0.665 ;
        RECT  2.260 0.530 2.370 1.140 ;
        RECT  1.910 1.035 2.260 1.140 ;
        RECT  1.800 0.885 1.910 1.140 ;
        RECT  1.710 0.480 1.835 0.595 ;
        RECT  1.710 1.230 1.760 1.475 ;
        RECT  1.620 0.480 1.710 1.475 ;
        RECT  1.440 0.390 1.530 1.395 ;
        RECT  1.405 0.390 1.440 0.595 ;
        RECT  0.945 1.305 1.440 1.395 ;
        RECT  0.830 0.495 1.405 0.595 ;
        RECT  0.695 0.295 1.295 0.405 ;
        RECT  0.560 0.865 1.140 0.975 ;
        RECT  0.840 1.305 0.945 1.495 ;
        RECT  0.585 0.295 0.695 0.505 ;
        RECT  0.440 0.865 0.560 1.195 ;
        RECT  0.350 0.865 0.440 0.965 ;
        RECT  0.260 0.500 0.350 1.385 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.275 0.260 1.385 ;
        RECT  0.075 0.285 0.185 0.590 ;
        RECT  0.075 1.275 0.185 1.465 ;
    END
END SDFKCSND2

MACRO SDFKCSND4
    CLASS CORE ;
    FOREIGN SDFKCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.500 2.150 0.930 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0539 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.275 2.755 0.690 ;
        RECT  2.415 0.275 2.635 0.440 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.745 0.295 8.875 0.675 ;
        RECT  8.745 1.020 8.875 1.470 ;
        RECT  8.650 0.525 8.745 0.675 ;
        RECT  8.650 1.020 8.745 1.190 ;
        RECT  8.355 0.525 8.650 1.190 ;
        RECT  8.350 0.295 8.355 1.490 ;
        RECT  8.225 0.295 8.350 0.675 ;
        RECT  8.225 1.020 8.350 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.945 7.875 1.115 ;
        RECT  7.705 0.295 7.835 0.710 ;
        RECT  7.650 0.540 7.705 0.710 ;
        RECT  7.350 0.540 7.650 1.115 ;
        RECT  7.315 0.540 7.350 0.710 ;
        RECT  7.145 0.945 7.350 1.115 ;
        RECT  7.185 0.295 7.315 0.710 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.065 0.880 1.175 ;
        RECT  0.650 1.065 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.710 3.345 0.890 ;
        RECT  2.895 0.710 2.995 1.290 ;
        RECT  2.845 1.060 2.895 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.685 1.350 1.215 ;
        RECT  0.630 0.685 1.250 0.775 ;
        RECT  0.990 1.105 1.250 1.215 ;
        RECT  0.460 0.660 0.630 0.775 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.135 -0.165 9.200 0.165 ;
        RECT  9.005 -0.165 9.135 0.695 ;
        RECT  8.635 -0.165 9.005 0.165 ;
        RECT  8.465 -0.165 8.635 0.425 ;
        RECT  8.095 -0.165 8.465 0.165 ;
        RECT  7.965 -0.165 8.095 0.675 ;
        RECT  7.575 -0.165 7.965 0.165 ;
        RECT  7.435 -0.165 7.575 0.450 ;
        RECT  6.550 -0.165 7.435 0.165 ;
        RECT  6.440 -0.165 6.550 0.450 ;
        RECT  5.275 -0.165 6.440 0.165 ;
        RECT  5.165 -0.165 5.275 0.625 ;
        RECT  4.660 -0.165 5.165 0.165 ;
        RECT  4.660 0.330 4.780 0.440 ;
        RECT  4.570 -0.165 4.660 0.440 ;
        RECT  2.270 -0.165 4.570 0.165 ;
        RECT  2.150 -0.165 2.270 0.395 ;
        RECT  0.000 -0.165 2.150 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.135 1.635 9.200 1.965 ;
        RECT  9.005 1.035 9.135 1.965 ;
        RECT  8.615 1.635 9.005 1.965 ;
        RECT  8.485 1.325 8.615 1.965 ;
        RECT  8.115 1.635 8.485 1.965 ;
        RECT  7.945 1.385 8.115 1.965 ;
        RECT  7.595 1.635 7.945 1.965 ;
        RECT  7.425 1.385 7.595 1.965 ;
        RECT  6.515 1.635 7.425 1.965 ;
        RECT  6.405 1.250 6.515 1.965 ;
        RECT  5.155 1.635 6.405 1.965 ;
        RECT  5.155 1.215 5.235 1.305 ;
        RECT  5.065 1.215 5.155 1.965 ;
        RECT  4.725 1.635 5.065 1.965 ;
        RECT  4.545 1.215 4.725 1.965 ;
        RECT  2.685 1.635 4.545 1.965 ;
        RECT  2.555 1.440 2.685 1.965 ;
        RECT  2.300 1.635 2.555 1.965 ;
        RECT  2.130 1.415 2.300 1.965 ;
        RECT  1.260 1.635 2.130 1.965 ;
        RECT  1.090 1.495 1.260 1.965 ;
        RECT  0.500 1.635 1.090 1.965 ;
        RECT  0.330 1.495 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.745 0.295 8.875 0.675 ;
        RECT  8.750 1.020 8.875 1.470 ;
        RECT  8.225 0.295 8.250 0.675 ;
        RECT  8.225 1.020 8.250 1.490 ;
        RECT  7.750 0.945 7.875 1.115 ;
        RECT  7.750 0.295 7.835 0.710 ;
        RECT  7.185 0.295 7.250 0.710 ;
        RECT  7.145 0.945 7.250 1.115 ;
        RECT  8.085 0.800 8.250 0.910 ;
        RECT  7.995 0.800 8.085 1.295 ;
        RECT  6.830 1.205 7.995 1.295 ;
        RECT  6.735 0.255 6.830 1.480 ;
        RECT  6.695 0.255 6.735 0.710 ;
        RECT  6.690 1.250 6.735 1.480 ;
        RECT  6.295 0.600 6.695 0.710 ;
        RECT  6.525 0.855 6.635 1.085 ;
        RECT  6.300 0.855 6.525 0.945 ;
        RECT  6.210 0.855 6.300 1.495 ;
        RECT  6.200 0.855 6.210 0.955 ;
        RECT  5.465 1.385 6.210 1.495 ;
        RECT  6.110 0.275 6.200 0.955 ;
        RECT  6.005 1.090 6.120 1.270 ;
        RECT  5.925 0.275 6.110 0.415 ;
        RECT  5.895 0.560 6.005 1.270 ;
        RECT  5.535 0.275 5.925 0.365 ;
        RECT  5.725 0.455 5.795 0.895 ;
        RECT  5.685 0.455 5.725 1.270 ;
        RECT  5.615 0.805 5.685 1.270 ;
        RECT  5.020 0.805 5.615 0.895 ;
        RECT  5.425 0.275 5.535 0.640 ;
        RECT  5.355 1.075 5.465 1.495 ;
        RECT  4.945 0.455 5.020 1.110 ;
        RECT  4.930 0.455 4.945 1.285 ;
        RECT  4.915 0.455 4.930 0.625 ;
        RECT  4.835 1.020 4.930 1.285 ;
        RECT  4.790 0.740 4.840 0.910 ;
        RECT  4.590 1.020 4.835 1.110 ;
        RECT  4.700 0.540 4.790 0.910 ;
        RECT  4.220 0.540 4.700 0.630 ;
        RECT  4.480 0.740 4.590 1.110 ;
        RECT  4.110 0.330 4.220 1.365 ;
        RECT  3.920 0.265 4.010 1.525 ;
        RECT  3.795 0.265 3.920 0.375 ;
        RECT  3.050 1.435 3.920 1.525 ;
        RECT  3.740 0.485 3.830 1.295 ;
        RECT  3.035 0.275 3.795 0.375 ;
        RECT  3.620 0.485 3.740 0.655 ;
        RECT  3.560 1.160 3.740 1.295 ;
        RECT  3.530 0.735 3.555 1.070 ;
        RECT  3.435 0.510 3.530 1.070 ;
        RECT  3.055 0.510 3.435 0.620 ;
        RECT  3.220 0.980 3.435 1.070 ;
        RECT  3.110 0.980 3.220 1.250 ;
        RECT  2.835 1.415 3.050 1.525 ;
        RECT  2.845 0.265 3.035 0.375 ;
        RECT  2.700 0.780 2.805 0.950 ;
        RECT  2.610 0.780 2.700 1.320 ;
        RECT  1.760 1.230 2.610 1.320 ;
        RECT  2.370 1.030 2.510 1.140 ;
        RECT  2.370 0.530 2.490 0.665 ;
        RECT  2.260 0.530 2.370 1.140 ;
        RECT  1.910 1.035 2.260 1.140 ;
        RECT  1.800 0.885 1.910 1.140 ;
        RECT  1.710 0.480 1.835 0.595 ;
        RECT  1.710 1.230 1.760 1.475 ;
        RECT  1.620 0.480 1.710 1.475 ;
        RECT  1.440 0.390 1.530 1.395 ;
        RECT  1.405 0.390 1.440 0.595 ;
        RECT  0.945 1.305 1.440 1.395 ;
        RECT  0.830 0.495 1.405 0.595 ;
        RECT  0.695 0.295 1.295 0.405 ;
        RECT  0.560 0.865 1.140 0.975 ;
        RECT  0.840 1.305 0.945 1.495 ;
        RECT  0.585 0.295 0.695 0.505 ;
        RECT  0.440 0.865 0.560 1.195 ;
        RECT  0.350 0.865 0.440 0.965 ;
        RECT  0.260 0.500 0.350 1.385 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.275 0.260 1.385 ;
        RECT  0.075 0.285 0.185 0.590 ;
        RECT  0.075 1.275 0.185 1.465 ;
    END
END SDFKCSND4

MACRO SDFKCSNQD0
    CLASS CORE ;
    FOREIGN SDFKCSNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.910 1.350 1.090 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.035 0.710 3.185 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0516 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.635 0.710 1.750 1.090 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0180 ;
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.460 0.400 6.550 1.525 ;
        RECT  6.415 0.400 6.460 0.640 ;
        RECT  6.410 1.040 6.460 1.525 ;
        RECT  6.130 0.550 6.415 0.640 ;
        RECT  6.020 0.550 6.130 0.955 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0342 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.710 0.600 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 0.710 3.570 1.090 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0342 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.720 0.290 0.830 ;
        RECT  0.045 0.310 0.170 0.830 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.275 -0.165 6.600 0.165 ;
        RECT  6.145 -0.165 6.275 0.445 ;
        RECT  2.125 -0.165 6.145 0.165 ;
        RECT  1.955 -0.165 2.125 0.405 ;
        RECT  0.000 -0.165 1.955 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.295 1.635 6.600 1.965 ;
        RECT  6.115 1.395 6.295 1.965 ;
        RECT  5.095 1.635 6.115 1.965 ;
        RECT  4.925 1.380 5.095 1.965 ;
        RECT  0.370 1.635 4.925 1.965 ;
        RECT  0.280 1.395 0.370 1.965 ;
        RECT  0.090 1.395 0.280 1.495 ;
        RECT  0.000 1.635 0.280 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.320 0.730 6.370 0.930 ;
        RECT  6.230 0.730 6.320 1.295 ;
        RECT  5.655 1.205 6.230 1.295 ;
        RECT  5.775 0.275 5.875 1.115 ;
        RECT  5.565 0.275 5.775 0.365 ;
        RECT  5.545 0.480 5.655 1.515 ;
        RECT  5.355 0.255 5.565 0.365 ;
        RECT  5.510 0.480 5.545 0.770 ;
        RECT  5.285 0.510 5.395 1.520 ;
        RECT  4.745 0.275 5.355 0.365 ;
        RECT  4.945 0.510 5.285 0.620 ;
        RECT  5.085 0.740 5.195 1.230 ;
        RECT  4.575 1.120 5.085 1.230 ;
        RECT  4.835 0.510 4.945 0.940 ;
        RECT  4.535 0.255 4.745 0.365 ;
        RECT  4.465 0.475 4.575 1.230 ;
        RECT  4.400 1.120 4.465 1.230 ;
        RECT  4.060 0.795 4.320 0.925 ;
        RECT  4.170 0.275 4.300 0.515 ;
        RECT  4.180 1.070 4.290 1.525 ;
        RECT  2.530 1.435 4.180 1.525 ;
        RECT  2.610 0.275 4.170 0.365 ;
        RECT  3.955 0.485 4.060 1.325 ;
        RECT  3.880 0.485 3.955 0.595 ;
        RECT  3.920 1.080 3.955 1.325 ;
        RECT  3.770 0.750 3.865 0.920 ;
        RECT  3.680 0.510 3.770 1.290 ;
        RECT  3.390 0.510 3.680 0.620 ;
        RECT  3.390 1.180 3.680 1.290 ;
        RECT  2.925 0.510 3.300 0.620 ;
        RECT  2.925 1.180 3.300 1.290 ;
        RECT  2.815 0.510 2.925 1.290 ;
        RECT  2.555 0.725 2.665 1.090 ;
        RECT  2.440 0.275 2.610 0.620 ;
        RECT  1.955 0.725 2.555 0.815 ;
        RECT  2.420 1.215 2.530 1.525 ;
        RECT  2.230 0.950 2.445 1.060 ;
        RECT  2.110 0.950 2.230 1.495 ;
        RECT  1.530 1.385 2.110 1.495 ;
        RECT  1.840 0.510 1.955 1.290 ;
        RECT  1.835 0.510 1.840 0.600 ;
        RECT  1.670 1.180 1.840 1.290 ;
        RECT  1.725 0.360 1.835 0.600 ;
        RECT  1.440 0.275 1.530 1.495 ;
        RECT  0.570 0.275 1.440 0.385 ;
        RECT  0.590 1.385 1.440 1.495 ;
        RECT  1.225 0.475 1.335 0.780 ;
        RECT  0.860 1.190 1.330 1.280 ;
        RECT  0.860 0.690 1.225 0.780 ;
        RECT  0.305 0.485 1.045 0.595 ;
        RECT  0.750 0.690 0.860 1.280 ;
        RECT  0.295 1.190 0.750 1.280 ;
        RECT  0.185 0.930 0.295 1.280 ;
    END
END SDFKCSNQD0

MACRO SDFKCSNQD1
    CLASS CORE ;
    FOREIGN SDFKCSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.500 2.150 0.930 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0539 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.275 2.755 0.690 ;
        RECT  2.415 0.275 2.635 0.440 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.255 0.560 6.355 1.110 ;
        RECT  6.245 0.280 6.255 1.440 ;
        RECT  6.145 0.280 6.245 0.685 ;
        RECT  6.145 0.985 6.245 1.440 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.065 0.880 1.175 ;
        RECT  0.650 1.065 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.710 3.320 0.890 ;
        RECT  2.895 0.710 2.995 1.290 ;
        RECT  2.845 1.060 2.895 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.685 1.350 1.215 ;
        RECT  0.630 0.685 1.250 0.775 ;
        RECT  0.990 1.105 1.250 1.215 ;
        RECT  0.460 0.660 0.630 0.775 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.515 -0.165 6.600 0.165 ;
        RECT  6.405 -0.165 6.515 0.445 ;
        RECT  5.720 -0.165 6.405 0.165 ;
        RECT  5.610 -0.165 5.720 0.450 ;
        RECT  4.610 -0.165 5.610 0.165 ;
        RECT  4.610 0.385 4.730 0.495 ;
        RECT  4.520 -0.165 4.610 0.495 ;
        RECT  2.270 -0.165 4.520 0.165 ;
        RECT  2.160 -0.165 2.270 0.395 ;
        RECT  0.000 -0.165 2.160 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.515 1.635 6.600 1.965 ;
        RECT  6.405 1.265 6.515 1.965 ;
        RECT  5.685 1.635 6.405 1.965 ;
        RECT  5.575 1.330 5.685 1.965 ;
        RECT  4.675 1.635 5.575 1.965 ;
        RECT  4.495 1.215 4.675 1.965 ;
        RECT  2.685 1.635 4.495 1.965 ;
        RECT  2.555 1.440 2.685 1.965 ;
        RECT  2.300 1.635 2.555 1.965 ;
        RECT  2.130 1.415 2.300 1.965 ;
        RECT  1.260 1.635 2.130 1.965 ;
        RECT  1.090 1.495 1.260 1.965 ;
        RECT  0.500 1.635 1.090 1.965 ;
        RECT  0.330 1.495 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.905 0.255 6.010 1.545 ;
        RECT  5.870 0.255 5.905 0.710 ;
        RECT  5.860 1.335 5.905 1.545 ;
        RECT  5.465 0.600 5.870 0.710 ;
        RECT  5.695 0.855 5.805 1.085 ;
        RECT  5.470 0.855 5.695 0.945 ;
        RECT  5.380 0.855 5.470 1.495 ;
        RECT  5.370 0.855 5.380 0.955 ;
        RECT  4.995 1.385 5.380 1.495 ;
        RECT  5.280 0.305 5.370 0.955 ;
        RECT  5.170 1.090 5.290 1.270 ;
        RECT  5.090 0.305 5.280 0.415 ;
        RECT  5.060 0.560 5.170 1.270 ;
        RECT  4.895 0.465 4.970 1.110 ;
        RECT  4.880 0.465 4.895 1.285 ;
        RECT  4.865 0.465 4.880 0.635 ;
        RECT  4.785 1.020 4.880 1.285 ;
        RECT  4.740 0.740 4.790 0.910 ;
        RECT  4.540 1.020 4.785 1.110 ;
        RECT  4.650 0.595 4.740 0.910 ;
        RECT  4.170 0.595 4.650 0.685 ;
        RECT  4.430 0.795 4.540 1.110 ;
        RECT  4.060 0.330 4.170 1.365 ;
        RECT  3.870 0.265 3.960 1.525 ;
        RECT  3.745 0.265 3.870 0.375 ;
        RECT  3.050 1.435 3.870 1.525 ;
        RECT  3.690 0.485 3.780 1.275 ;
        RECT  3.035 0.275 3.745 0.375 ;
        RECT  3.595 0.485 3.690 0.655 ;
        RECT  3.535 1.165 3.690 1.275 ;
        RECT  3.505 0.735 3.530 1.070 ;
        RECT  3.410 0.510 3.505 1.070 ;
        RECT  3.055 0.510 3.410 0.620 ;
        RECT  3.195 0.980 3.410 1.070 ;
        RECT  3.085 0.980 3.195 1.250 ;
        RECT  2.835 1.415 3.050 1.525 ;
        RECT  2.845 0.265 3.035 0.375 ;
        RECT  2.700 0.780 2.805 0.950 ;
        RECT  2.610 0.780 2.700 1.320 ;
        RECT  1.750 1.230 2.610 1.320 ;
        RECT  2.370 1.030 2.510 1.140 ;
        RECT  2.370 0.545 2.490 0.655 ;
        RECT  2.260 0.545 2.370 1.140 ;
        RECT  1.910 1.035 2.260 1.140 ;
        RECT  1.800 0.885 1.910 1.140 ;
        RECT  1.710 0.485 1.835 0.595 ;
        RECT  1.710 1.230 1.750 1.475 ;
        RECT  1.620 0.485 1.710 1.475 ;
        RECT  1.440 0.390 1.530 1.395 ;
        RECT  1.405 0.390 1.440 0.595 ;
        RECT  0.945 1.305 1.440 1.395 ;
        RECT  0.830 0.495 1.405 0.595 ;
        RECT  0.695 0.295 1.295 0.405 ;
        RECT  0.560 0.865 1.140 0.975 ;
        RECT  0.840 1.305 0.945 1.495 ;
        RECT  0.585 0.295 0.695 0.505 ;
        RECT  0.440 0.865 0.560 1.195 ;
        RECT  0.350 0.865 0.440 0.965 ;
        RECT  0.260 0.500 0.350 1.385 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.275 0.260 1.385 ;
        RECT  0.075 0.280 0.185 0.590 ;
        RECT  0.075 1.275 0.185 1.465 ;
    END
END SDFKCSNQD1

MACRO SDFKCSNQD2
    CLASS CORE ;
    FOREIGN SDFKCSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.500 2.150 0.930 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0539 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.275 2.755 0.690 ;
        RECT  2.415 0.275 2.635 0.440 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.355 0.285 6.465 0.700 ;
        RECT  6.355 1.045 6.465 1.460 ;
        RECT  6.250 0.545 6.355 1.165 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.065 0.880 1.175 ;
        RECT  0.650 1.065 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.710 3.320 0.890 ;
        RECT  2.895 0.710 2.995 1.290 ;
        RECT  2.845 1.060 2.895 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.685 1.350 1.215 ;
        RECT  0.630 0.685 1.250 0.775 ;
        RECT  0.990 1.105 1.250 1.215 ;
        RECT  0.460 0.660 0.630 0.775 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 -0.165 6.800 0.165 ;
        RECT  6.615 -0.165 6.725 0.675 ;
        RECT  5.720 -0.165 6.615 0.165 ;
        RECT  5.610 -0.165 5.720 0.450 ;
        RECT  4.610 -0.165 5.610 0.165 ;
        RECT  4.610 0.385 4.730 0.495 ;
        RECT  4.520 -0.165 4.610 0.495 ;
        RECT  2.270 -0.165 4.520 0.165 ;
        RECT  2.150 -0.165 2.270 0.395 ;
        RECT  0.000 -0.165 2.150 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.725 1.635 6.800 1.965 ;
        RECT  6.615 1.045 6.725 1.965 ;
        RECT  5.685 1.635 6.615 1.965 ;
        RECT  5.575 1.330 5.685 1.965 ;
        RECT  4.675 1.635 5.575 1.965 ;
        RECT  4.495 1.215 4.675 1.965 ;
        RECT  2.685 1.635 4.495 1.965 ;
        RECT  2.555 1.440 2.685 1.965 ;
        RECT  2.300 1.635 2.555 1.965 ;
        RECT  2.130 1.415 2.300 1.965 ;
        RECT  1.260 1.635 2.130 1.965 ;
        RECT  1.090 1.495 1.260 1.965 ;
        RECT  0.500 1.635 1.090 1.965 ;
        RECT  0.330 1.495 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.905 0.255 6.015 1.545 ;
        RECT  5.870 0.255 5.905 0.710 ;
        RECT  5.860 1.315 5.905 1.545 ;
        RECT  5.465 0.600 5.870 0.710 ;
        RECT  5.695 0.855 5.805 1.085 ;
        RECT  5.470 0.855 5.695 0.945 ;
        RECT  5.380 0.855 5.470 1.495 ;
        RECT  5.370 0.855 5.380 0.955 ;
        RECT  4.995 1.380 5.380 1.495 ;
        RECT  5.280 0.305 5.370 0.955 ;
        RECT  5.170 1.090 5.290 1.270 ;
        RECT  5.090 0.305 5.280 0.415 ;
        RECT  5.060 0.560 5.170 1.270 ;
        RECT  4.895 0.465 4.970 1.110 ;
        RECT  4.880 0.465 4.895 1.285 ;
        RECT  4.865 0.465 4.880 0.635 ;
        RECT  4.785 1.020 4.880 1.285 ;
        RECT  4.740 0.740 4.790 0.910 ;
        RECT  4.540 1.020 4.785 1.110 ;
        RECT  4.650 0.595 4.740 0.910 ;
        RECT  4.170 0.595 4.650 0.685 ;
        RECT  4.430 0.795 4.540 1.110 ;
        RECT  4.060 0.330 4.170 1.365 ;
        RECT  3.870 0.265 3.960 1.525 ;
        RECT  3.745 0.265 3.870 0.375 ;
        RECT  3.050 1.435 3.870 1.525 ;
        RECT  3.690 0.485 3.780 1.295 ;
        RECT  3.035 0.275 3.745 0.375 ;
        RECT  3.595 0.485 3.690 0.655 ;
        RECT  3.535 1.160 3.690 1.295 ;
        RECT  3.505 0.735 3.530 1.070 ;
        RECT  3.410 0.510 3.505 1.070 ;
        RECT  3.055 0.510 3.410 0.620 ;
        RECT  3.195 0.980 3.410 1.070 ;
        RECT  3.085 0.980 3.195 1.250 ;
        RECT  2.835 1.415 3.050 1.525 ;
        RECT  2.845 0.265 3.035 0.375 ;
        RECT  2.700 0.780 2.805 0.950 ;
        RECT  2.610 0.780 2.700 1.320 ;
        RECT  1.760 1.230 2.610 1.320 ;
        RECT  2.370 1.030 2.510 1.140 ;
        RECT  2.370 0.530 2.490 0.665 ;
        RECT  2.260 0.530 2.370 1.140 ;
        RECT  1.910 1.035 2.260 1.140 ;
        RECT  1.800 0.885 1.910 1.140 ;
        RECT  1.710 0.480 1.835 0.595 ;
        RECT  1.710 1.230 1.760 1.475 ;
        RECT  1.620 0.480 1.710 1.475 ;
        RECT  1.440 0.390 1.530 1.395 ;
        RECT  1.405 0.390 1.440 0.595 ;
        RECT  0.945 1.305 1.440 1.395 ;
        RECT  0.830 0.495 1.405 0.595 ;
        RECT  0.695 0.295 1.295 0.405 ;
        RECT  0.560 0.865 1.140 0.975 ;
        RECT  0.840 1.305 0.945 1.495 ;
        RECT  0.585 0.295 0.695 0.505 ;
        RECT  0.440 0.865 0.560 1.195 ;
        RECT  0.350 0.865 0.440 0.965 ;
        RECT  0.260 0.500 0.350 1.385 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.275 0.260 1.385 ;
        RECT  0.075 0.285 0.185 0.590 ;
        RECT  0.075 1.275 0.185 1.465 ;
    END
END SDFKCSNQD2

MACRO SDFKCSNQD4
    CLASS CORE ;
    FOREIGN SDFKCSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.500 2.150 0.930 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0539 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.275 2.755 0.690 ;
        RECT  2.415 0.275 2.635 0.440 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.755 0.295 7.865 0.675 ;
        RECT  7.755 1.020 7.865 1.460 ;
        RECT  7.650 0.525 7.755 0.675 ;
        RECT  7.650 1.020 7.755 1.190 ;
        RECT  7.350 0.525 7.650 1.190 ;
        RECT  7.345 0.525 7.350 0.675 ;
        RECT  7.345 1.020 7.350 1.190 ;
        RECT  7.235 0.295 7.345 0.675 ;
        RECT  7.235 1.020 7.345 1.460 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0286 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.065 0.880 1.175 ;
        RECT  0.650 1.065 0.750 1.500 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.710 3.345 0.890 ;
        RECT  2.895 0.710 2.995 1.290 ;
        RECT  2.845 1.060 2.895 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.685 1.350 1.215 ;
        RECT  0.630 0.685 1.250 0.775 ;
        RECT  0.990 1.105 1.250 1.215 ;
        RECT  0.460 0.660 0.630 0.775 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.125 -0.165 8.200 0.165 ;
        RECT  8.015 -0.165 8.125 0.695 ;
        RECT  7.635 -0.165 8.015 0.165 ;
        RECT  7.465 -0.165 7.635 0.425 ;
        RECT  7.085 -0.165 7.465 0.165 ;
        RECT  6.975 -0.165 7.085 0.680 ;
        RECT  6.550 -0.165 6.975 0.165 ;
        RECT  6.440 -0.165 6.550 0.450 ;
        RECT  5.275 -0.165 6.440 0.165 ;
        RECT  5.165 -0.165 5.275 0.625 ;
        RECT  4.660 -0.165 5.165 0.165 ;
        RECT  4.660 0.330 4.780 0.440 ;
        RECT  4.570 -0.165 4.660 0.440 ;
        RECT  2.270 -0.165 4.570 0.165 ;
        RECT  2.150 -0.165 2.270 0.395 ;
        RECT  0.000 -0.165 2.150 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.125 1.635 8.200 1.965 ;
        RECT  8.015 1.050 8.125 1.965 ;
        RECT  7.605 1.635 8.015 1.965 ;
        RECT  7.495 1.325 7.605 1.965 ;
        RECT  7.085 1.635 7.495 1.965 ;
        RECT  6.975 1.045 7.085 1.965 ;
        RECT  6.515 1.635 6.975 1.965 ;
        RECT  6.405 1.330 6.515 1.965 ;
        RECT  5.155 1.635 6.405 1.965 ;
        RECT  5.155 1.215 5.235 1.305 ;
        RECT  5.065 1.215 5.155 1.965 ;
        RECT  4.725 1.635 5.065 1.965 ;
        RECT  4.545 1.215 4.725 1.965 ;
        RECT  2.685 1.635 4.545 1.965 ;
        RECT  2.555 1.440 2.685 1.965 ;
        RECT  2.300 1.635 2.555 1.965 ;
        RECT  2.130 1.415 2.300 1.965 ;
        RECT  1.260 1.635 2.130 1.965 ;
        RECT  1.090 1.495 1.260 1.965 ;
        RECT  0.500 1.635 1.090 1.965 ;
        RECT  0.330 1.495 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.755 0.295 7.865 0.675 ;
        RECT  7.755 1.020 7.865 1.460 ;
        RECT  7.750 0.525 7.755 0.675 ;
        RECT  7.750 1.020 7.755 1.190 ;
        RECT  7.235 0.295 7.250 0.675 ;
        RECT  7.235 1.020 7.250 1.460 ;
        RECT  6.735 0.255 6.850 1.545 ;
        RECT  6.700 0.255 6.735 0.710 ;
        RECT  6.690 1.315 6.735 1.545 ;
        RECT  6.295 0.600 6.700 0.710 ;
        RECT  6.525 0.855 6.635 1.085 ;
        RECT  6.300 0.855 6.525 0.945 ;
        RECT  6.210 0.855 6.300 1.495 ;
        RECT  6.200 0.855 6.210 0.955 ;
        RECT  5.465 1.385 6.210 1.495 ;
        RECT  6.110 0.275 6.200 0.955 ;
        RECT  6.005 1.090 6.120 1.270 ;
        RECT  5.925 0.275 6.110 0.415 ;
        RECT  5.895 0.560 6.005 1.270 ;
        RECT  5.535 0.275 5.925 0.365 ;
        RECT  5.725 0.455 5.795 0.895 ;
        RECT  5.685 0.455 5.725 1.270 ;
        RECT  5.615 0.805 5.685 1.270 ;
        RECT  5.020 0.805 5.615 0.895 ;
        RECT  5.425 0.275 5.535 0.640 ;
        RECT  5.355 1.075 5.465 1.495 ;
        RECT  4.945 0.455 5.020 1.110 ;
        RECT  4.930 0.455 4.945 1.285 ;
        RECT  4.915 0.455 4.930 0.625 ;
        RECT  4.835 1.020 4.930 1.285 ;
        RECT  4.790 0.740 4.840 0.910 ;
        RECT  4.590 1.020 4.835 1.110 ;
        RECT  4.700 0.540 4.790 0.910 ;
        RECT  4.220 0.540 4.700 0.630 ;
        RECT  4.480 0.740 4.590 1.110 ;
        RECT  4.110 0.330 4.220 1.365 ;
        RECT  3.920 0.265 4.010 1.525 ;
        RECT  3.795 0.265 3.920 0.375 ;
        RECT  3.050 1.435 3.920 1.525 ;
        RECT  3.740 0.485 3.830 1.295 ;
        RECT  3.035 0.275 3.795 0.375 ;
        RECT  3.620 0.485 3.740 0.655 ;
        RECT  3.560 1.160 3.740 1.295 ;
        RECT  3.530 0.735 3.555 1.070 ;
        RECT  3.435 0.510 3.530 1.070 ;
        RECT  3.055 0.510 3.435 0.620 ;
        RECT  3.220 0.980 3.435 1.070 ;
        RECT  3.110 0.980 3.220 1.250 ;
        RECT  2.835 1.415 3.050 1.525 ;
        RECT  2.845 0.265 3.035 0.375 ;
        RECT  2.700 0.780 2.805 0.950 ;
        RECT  2.610 0.780 2.700 1.320 ;
        RECT  1.760 1.230 2.610 1.320 ;
        RECT  2.370 1.030 2.510 1.140 ;
        RECT  2.370 0.530 2.490 0.665 ;
        RECT  2.260 0.530 2.370 1.140 ;
        RECT  1.910 1.035 2.260 1.140 ;
        RECT  1.800 0.885 1.910 1.140 ;
        RECT  1.710 0.480 1.835 0.595 ;
        RECT  1.710 1.230 1.760 1.475 ;
        RECT  1.620 0.480 1.710 1.475 ;
        RECT  1.440 0.390 1.530 1.395 ;
        RECT  1.405 0.390 1.440 0.595 ;
        RECT  0.945 1.305 1.440 1.395 ;
        RECT  0.830 0.495 1.405 0.595 ;
        RECT  0.695 0.295 1.295 0.405 ;
        RECT  0.560 0.865 1.140 0.975 ;
        RECT  0.840 1.305 0.945 1.495 ;
        RECT  0.585 0.295 0.695 0.505 ;
        RECT  0.440 0.865 0.560 1.195 ;
        RECT  0.350 0.865 0.440 0.965 ;
        RECT  0.260 0.500 0.350 1.385 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.275 0.260 1.385 ;
        RECT  0.075 0.285 0.185 0.590 ;
        RECT  0.075 1.275 0.185 1.465 ;
    END
END SDFKCSNQD4

MACRO SDFKSND0
    CLASS CORE ;
    FOREIGN SDFKSND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.775 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0539 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.310 2.350 0.690 ;
        RECT  2.040 0.310 2.250 0.420 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.480 6.350 1.290 ;
        RECT  6.215 0.480 6.250 0.675 ;
        RECT  6.225 1.040 6.250 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.525 5.950 1.180 ;
        RECT  5.680 0.525 5.850 0.635 ;
        RECT  5.685 1.070 5.850 1.180 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.780 0.880 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 0.710 2.925 0.890 ;
        RECT  2.510 0.710 2.600 1.290 ;
        RECT  2.450 1.060 2.510 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 -0.165 6.400 0.165 ;
        RECT  4.175 -0.165 4.285 0.490 ;
        RECT  1.895 -0.165 4.175 0.165 ;
        RECT  1.785 -0.165 1.895 0.400 ;
        RECT  0.000 -0.165 1.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.290 1.635 6.400 1.965 ;
        RECT  5.180 1.250 5.290 1.965 ;
        RECT  4.280 1.635 5.180 1.965 ;
        RECT  4.100 1.200 4.280 1.965 ;
        RECT  2.300 1.635 4.100 1.965 ;
        RECT  2.190 1.440 2.300 1.965 ;
        RECT  1.730 1.635 2.190 1.965 ;
        RECT  1.560 1.395 1.730 1.965 ;
        RECT  0.475 1.635 1.560 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.135 0.775 6.160 0.945 ;
        RECT  6.045 0.775 6.135 1.390 ;
        RECT  5.590 1.290 6.045 1.390 ;
        RECT  5.575 0.600 5.590 1.390 ;
        RECT  5.565 0.600 5.575 1.545 ;
        RECT  5.500 0.265 5.565 1.545 ;
        RECT  5.455 0.265 5.500 0.710 ;
        RECT  5.465 1.290 5.500 1.545 ;
        RECT  5.070 0.600 5.455 0.710 ;
        RECT  5.300 0.855 5.410 1.085 ;
        RECT  5.085 0.855 5.300 0.945 ;
        RECT  4.995 0.855 5.085 1.495 ;
        RECT  4.975 0.855 4.995 0.945 ;
        RECT  4.600 1.380 4.995 1.495 ;
        RECT  4.885 0.305 4.975 0.945 ;
        RECT  4.780 1.090 4.905 1.260 ;
        RECT  4.695 0.305 4.885 0.415 ;
        RECT  4.670 0.565 4.780 1.260 ;
        RECT  4.500 0.465 4.575 1.110 ;
        RECT  4.485 0.465 4.500 1.285 ;
        RECT  4.460 0.465 4.485 0.635 ;
        RECT  4.390 1.020 4.485 1.285 ;
        RECT  4.345 0.740 4.395 0.910 ;
        RECT  4.145 1.020 4.390 1.110 ;
        RECT  4.255 0.590 4.345 0.910 ;
        RECT  3.775 0.590 4.255 0.680 ;
        RECT  4.035 0.785 4.145 1.110 ;
        RECT  3.665 0.330 3.775 1.365 ;
        RECT  3.475 0.255 3.565 1.525 ;
        RECT  3.350 0.255 3.475 0.375 ;
        RECT  2.480 1.415 3.475 1.525 ;
        RECT  3.275 0.485 3.385 1.275 ;
        RECT  2.660 0.275 3.350 0.375 ;
        RECT  3.200 0.485 3.275 0.655 ;
        RECT  3.140 1.165 3.275 1.275 ;
        RECT  3.110 0.735 3.145 0.905 ;
        RECT  3.015 0.515 3.110 1.070 ;
        RECT  2.650 0.515 3.015 0.620 ;
        RECT  2.800 0.980 3.015 1.070 ;
        RECT  2.690 0.980 2.800 1.250 ;
        RECT  2.490 0.265 2.660 0.375 ;
        RECT  2.325 0.785 2.420 0.955 ;
        RECT  2.235 0.785 2.325 1.305 ;
        RECT  1.145 1.215 2.235 1.305 ;
        RECT  2.085 1.015 2.135 1.125 ;
        RECT  1.975 0.515 2.085 1.125 ;
        RECT  1.345 1.035 1.975 1.125 ;
        RECT  1.310 0.455 1.420 0.795 ;
        RECT  1.235 0.905 1.345 1.125 ;
        RECT  1.145 0.705 1.310 0.795 ;
        RECT  0.960 0.475 1.210 0.585 ;
        RECT  1.055 0.705 1.145 1.365 ;
        RECT  0.895 0.375 0.960 1.290 ;
        RECT  0.870 0.375 0.895 1.520 ;
        RECT  0.525 0.375 0.870 0.485 ;
        RECT  0.785 1.200 0.870 1.520 ;
        RECT  0.350 0.750 0.530 0.920 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.075 0.350 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.520 ;
    END
END SDFKSND0

MACRO SDFKSND1
    CLASS CORE ;
    FOREIGN SDFKSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.775 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0604 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.290 2.350 0.690 ;
        RECT  2.060 0.290 2.250 0.400 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.285 6.350 1.490 ;
        RECT  6.215 0.285 6.250 0.675 ;
        RECT  6.220 1.050 6.250 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.565 5.950 1.210 ;
        RECT  5.825 0.565 5.850 0.675 ;
        RECT  5.675 1.100 5.850 1.210 ;
        RECT  5.715 0.285 5.825 0.675 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.780 0.925 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.610 0.710 2.925 0.890 ;
        RECT  2.520 0.710 2.610 1.290 ;
        RECT  2.450 1.060 2.520 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 -0.165 6.400 0.165 ;
        RECT  4.175 -0.165 4.285 0.490 ;
        RECT  1.895 -0.165 4.175 0.165 ;
        RECT  1.785 -0.165 1.895 0.400 ;
        RECT  0.000 -0.165 1.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.285 1.635 6.400 1.965 ;
        RECT  5.175 1.250 5.285 1.965 ;
        RECT  4.280 1.635 5.175 1.965 ;
        RECT  4.100 1.200 4.280 1.965 ;
        RECT  2.300 1.635 4.100 1.965 ;
        RECT  2.190 1.440 2.300 1.965 ;
        RECT  1.725 1.635 2.190 1.965 ;
        RECT  1.555 1.405 1.725 1.965 ;
        RECT  0.475 1.635 1.555 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.130 0.775 6.160 0.945 ;
        RECT  6.040 0.775 6.130 1.415 ;
        RECT  5.565 1.305 6.040 1.415 ;
        RECT  5.475 0.265 5.565 1.415 ;
        RECT  5.455 0.265 5.475 0.690 ;
        RECT  5.385 1.305 5.475 1.415 ;
        RECT  5.070 0.580 5.455 0.690 ;
        RECT  5.085 0.840 5.380 1.010 ;
        RECT  4.995 0.840 5.085 1.495 ;
        RECT  4.975 0.840 4.995 0.945 ;
        RECT  4.600 1.380 4.995 1.495 ;
        RECT  4.885 0.305 4.975 0.945 ;
        RECT  4.780 1.090 4.905 1.260 ;
        RECT  4.695 0.305 4.885 0.415 ;
        RECT  4.670 0.565 4.780 1.260 ;
        RECT  4.500 0.465 4.575 1.110 ;
        RECT  4.485 0.465 4.500 1.285 ;
        RECT  4.460 0.465 4.485 0.635 ;
        RECT  4.390 1.020 4.485 1.285 ;
        RECT  4.345 0.740 4.395 0.910 ;
        RECT  4.145 1.020 4.390 1.110 ;
        RECT  4.255 0.590 4.345 0.910 ;
        RECT  3.775 0.590 4.255 0.680 ;
        RECT  4.035 0.785 4.145 1.110 ;
        RECT  3.665 0.330 3.775 1.365 ;
        RECT  3.475 0.255 3.565 1.525 ;
        RECT  3.350 0.255 3.475 0.375 ;
        RECT  2.480 1.415 3.475 1.525 ;
        RECT  3.275 0.485 3.385 1.275 ;
        RECT  2.680 0.275 3.350 0.375 ;
        RECT  3.210 0.485 3.275 0.655 ;
        RECT  3.140 1.165 3.275 1.275 ;
        RECT  3.110 0.735 3.155 0.905 ;
        RECT  3.015 0.515 3.110 1.070 ;
        RECT  2.670 0.515 3.015 0.620 ;
        RECT  2.800 0.980 3.015 1.070 ;
        RECT  2.700 0.980 2.800 1.250 ;
        RECT  2.510 0.265 2.680 0.375 ;
        RECT  2.325 0.785 2.430 0.955 ;
        RECT  2.235 0.785 2.325 1.315 ;
        RECT  1.140 1.215 2.235 1.315 ;
        RECT  2.105 1.015 2.135 1.125 ;
        RECT  1.995 0.515 2.105 1.125 ;
        RECT  1.345 1.035 1.995 1.125 ;
        RECT  1.310 0.455 1.420 0.795 ;
        RECT  1.235 0.905 1.345 1.125 ;
        RECT  1.140 0.705 1.310 0.795 ;
        RECT  0.960 0.475 1.210 0.585 ;
        RECT  1.050 0.705 1.140 1.315 ;
        RECT  0.930 0.375 0.960 1.290 ;
        RECT  0.870 0.375 0.930 1.520 ;
        RECT  0.525 0.375 0.870 0.485 ;
        RECT  0.820 1.200 0.870 1.520 ;
        RECT  0.350 0.750 0.530 0.920 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.075 0.350 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.520 ;
    END
END SDFKSND1

MACRO SDFKSND2
    CLASS CORE ;
    FOREIGN SDFKSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.775 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0604 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.290 2.350 0.690 ;
        RECT  2.060 0.290 2.250 0.400 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.575 6.750 1.150 ;
        RECT  6.645 0.575 6.650 0.675 ;
        RECT  6.645 1.050 6.650 1.150 ;
        RECT  6.535 0.285 6.645 0.675 ;
        RECT  6.535 1.050 6.645 1.460 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.285 6.150 1.215 ;
        RECT  6.015 0.285 6.050 0.675 ;
        RECT  6.015 1.005 6.050 1.215 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.780 0.925 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.610 0.710 2.925 0.890 ;
        RECT  2.520 0.710 2.610 1.290 ;
        RECT  2.450 1.060 2.520 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.905 -0.165 7.000 0.165 ;
        RECT  6.795 -0.165 6.905 0.485 ;
        RECT  6.385 -0.165 6.795 0.165 ;
        RECT  6.275 -0.165 6.385 0.685 ;
        RECT  5.865 -0.165 6.275 0.165 ;
        RECT  5.755 -0.165 5.865 0.685 ;
        RECT  4.285 -0.165 5.755 0.165 ;
        RECT  4.175 -0.165 4.285 0.490 ;
        RECT  1.895 -0.165 4.175 0.165 ;
        RECT  1.785 -0.165 1.895 0.400 ;
        RECT  0.000 -0.165 1.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.905 1.635 7.000 1.965 ;
        RECT  6.795 1.250 6.905 1.965 ;
        RECT  5.870 1.635 6.795 1.965 ;
        RECT  5.700 1.505 5.870 1.965 ;
        RECT  5.285 1.635 5.700 1.965 ;
        RECT  5.175 1.250 5.285 1.965 ;
        RECT  4.280 1.635 5.175 1.965 ;
        RECT  4.100 1.200 4.280 1.965 ;
        RECT  2.300 1.635 4.100 1.965 ;
        RECT  2.190 1.440 2.300 1.965 ;
        RECT  1.725 1.635 2.190 1.965 ;
        RECT  1.555 1.405 1.725 1.965 ;
        RECT  0.475 1.635 1.555 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.425 0.805 6.540 0.915 ;
        RECT  6.335 0.805 6.425 1.415 ;
        RECT  5.565 1.305 6.335 1.415 ;
        RECT  5.475 0.265 5.565 1.415 ;
        RECT  5.455 0.265 5.475 0.690 ;
        RECT  5.385 1.305 5.475 1.415 ;
        RECT  5.070 0.580 5.455 0.690 ;
        RECT  5.085 0.840 5.380 1.010 ;
        RECT  4.995 0.840 5.085 1.495 ;
        RECT  4.975 0.840 4.995 0.945 ;
        RECT  4.600 1.380 4.995 1.495 ;
        RECT  4.885 0.305 4.975 0.945 ;
        RECT  4.780 1.090 4.905 1.260 ;
        RECT  4.695 0.305 4.885 0.415 ;
        RECT  4.670 0.565 4.780 1.260 ;
        RECT  4.500 0.465 4.575 1.110 ;
        RECT  4.485 0.465 4.500 1.285 ;
        RECT  4.460 0.465 4.485 0.635 ;
        RECT  4.390 1.020 4.485 1.285 ;
        RECT  4.345 0.740 4.395 0.910 ;
        RECT  4.145 1.020 4.390 1.110 ;
        RECT  4.255 0.590 4.345 0.910 ;
        RECT  3.775 0.590 4.255 0.680 ;
        RECT  4.035 0.785 4.145 1.110 ;
        RECT  3.665 0.330 3.775 1.365 ;
        RECT  3.475 0.255 3.565 1.525 ;
        RECT  3.350 0.255 3.475 0.375 ;
        RECT  2.480 1.415 3.475 1.525 ;
        RECT  3.275 0.485 3.385 1.275 ;
        RECT  2.680 0.275 3.350 0.375 ;
        RECT  3.210 0.485 3.275 0.655 ;
        RECT  3.140 1.165 3.275 1.275 ;
        RECT  3.110 0.735 3.155 0.905 ;
        RECT  3.015 0.515 3.110 1.070 ;
        RECT  2.670 0.515 3.015 0.620 ;
        RECT  2.800 0.980 3.015 1.070 ;
        RECT  2.700 0.980 2.800 1.250 ;
        RECT  2.510 0.265 2.680 0.375 ;
        RECT  2.325 0.785 2.430 0.955 ;
        RECT  2.235 0.785 2.325 1.315 ;
        RECT  1.140 1.215 2.235 1.315 ;
        RECT  2.105 1.015 2.135 1.125 ;
        RECT  1.995 0.515 2.105 1.125 ;
        RECT  1.345 1.035 1.995 1.125 ;
        RECT  1.310 0.455 1.420 0.795 ;
        RECT  1.235 0.905 1.345 1.125 ;
        RECT  1.140 0.705 1.310 0.795 ;
        RECT  0.960 0.475 1.210 0.585 ;
        RECT  1.050 0.705 1.140 1.315 ;
        RECT  0.930 0.375 0.960 1.290 ;
        RECT  0.870 0.375 0.930 1.520 ;
        RECT  0.525 0.375 0.870 0.485 ;
        RECT  0.820 1.200 0.870 1.520 ;
        RECT  0.350 0.750 0.530 0.920 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.075 0.350 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.520 ;
    END
END SDFKSND2

MACRO SDFKSND4
    CLASS CORE ;
    FOREIGN SDFKSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.775 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0604 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.290 2.350 0.690 ;
        RECT  2.060 0.290 2.250 0.400 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.355 0.295 8.465 0.675 ;
        RECT  8.355 1.020 8.465 1.470 ;
        RECT  8.250 0.525 8.355 0.675 ;
        RECT  8.250 1.020 8.355 1.190 ;
        RECT  7.950 0.525 8.250 1.190 ;
        RECT  7.945 0.525 7.950 0.675 ;
        RECT  7.835 1.020 7.950 1.490 ;
        RECT  7.835 0.295 7.945 0.675 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 1.070 7.485 1.240 ;
        RECT  7.250 0.325 7.475 0.645 ;
        RECT  6.950 0.325 7.250 1.240 ;
        RECT  6.785 0.325 6.950 0.645 ;
        RECT  6.775 1.070 6.950 1.240 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.780 0.925 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.815 0.510 2.950 0.910 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.725 -0.165 8.800 0.165 ;
        RECT  8.615 -0.165 8.725 0.695 ;
        RECT  8.235 -0.165 8.615 0.165 ;
        RECT  8.065 -0.165 8.235 0.435 ;
        RECT  4.940 -0.165 8.065 0.165 ;
        RECT  4.830 -0.165 4.940 0.685 ;
        RECT  4.325 -0.165 4.830 0.165 ;
        RECT  4.325 0.365 4.445 0.475 ;
        RECT  4.235 -0.165 4.325 0.475 ;
        RECT  1.895 -0.165 4.235 0.165 ;
        RECT  1.785 -0.165 1.895 0.400 ;
        RECT  0.000 -0.165 1.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.725 1.635 8.800 1.965 ;
        RECT  8.615 1.105 8.725 1.965 ;
        RECT  8.230 1.635 8.615 1.965 ;
        RECT  8.070 1.300 8.230 1.965 ;
        RECT  6.200 1.635 8.070 1.965 ;
        RECT  6.085 1.330 6.200 1.965 ;
        RECT  4.920 1.635 6.085 1.965 ;
        RECT  4.750 1.215 4.920 1.965 ;
        RECT  4.410 1.635 4.750 1.965 ;
        RECT  4.230 1.215 4.410 1.965 ;
        RECT  2.300 1.635 4.230 1.965 ;
        RECT  2.190 1.440 2.300 1.965 ;
        RECT  1.725 1.635 2.190 1.965 ;
        RECT  1.555 1.405 1.725 1.965 ;
        RECT  0.475 1.635 1.555 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.355 0.295 8.465 0.675 ;
        RECT  8.355 1.020 8.465 1.470 ;
        RECT  8.350 0.525 8.355 0.675 ;
        RECT  8.350 1.020 8.355 1.190 ;
        RECT  7.835 0.295 7.850 0.675 ;
        RECT  7.835 1.020 7.850 1.490 ;
        RECT  7.350 1.070 7.485 1.240 ;
        RECT  7.350 0.325 7.475 0.645 ;
        RECT  6.785 0.325 6.850 0.645 ;
        RECT  6.775 1.070 6.850 1.240 ;
        RECT  7.685 0.800 7.850 0.910 ;
        RECT  7.595 0.800 7.685 1.455 ;
        RECT  6.630 1.365 7.595 1.455 ;
        RECT  6.525 0.635 6.630 1.455 ;
        RECT  6.460 0.635 6.525 0.745 ;
        RECT  6.300 1.345 6.525 1.455 ;
        RECT  6.350 0.340 6.460 0.745 ;
        RECT  5.995 0.855 6.415 0.965 ;
        RECT  5.970 0.635 6.350 0.745 ;
        RECT  5.905 0.855 5.995 1.495 ;
        RECT  5.870 0.855 5.905 0.955 ;
        RECT  5.150 1.385 5.905 1.495 ;
        RECT  5.780 0.275 5.870 0.955 ;
        RECT  5.705 1.090 5.815 1.270 ;
        RECT  5.600 0.275 5.780 0.415 ;
        RECT  5.685 1.090 5.705 1.180 ;
        RECT  5.575 0.560 5.685 1.180 ;
        RECT  5.190 0.275 5.600 0.365 ;
        RECT  5.410 0.455 5.475 0.625 ;
        RECT  5.320 0.455 5.410 1.270 ;
        RECT  5.300 0.790 5.320 1.270 ;
        RECT  4.705 0.790 5.300 0.880 ;
        RECT  5.080 0.275 5.190 0.465 ;
        RECT  5.040 1.045 5.150 1.495 ;
        RECT  4.630 0.465 4.705 1.110 ;
        RECT  4.615 0.465 4.630 1.285 ;
        RECT  4.570 0.465 4.615 0.635 ;
        RECT  4.520 1.020 4.615 1.285 ;
        RECT  4.445 0.740 4.525 0.910 ;
        RECT  4.265 1.020 4.520 1.110 ;
        RECT  4.355 0.575 4.445 0.910 ;
        RECT  3.885 0.575 4.355 0.665 ;
        RECT  4.165 0.775 4.265 1.110 ;
        RECT  3.775 0.325 3.885 1.365 ;
        RECT  3.565 0.315 3.655 1.470 ;
        RECT  3.515 0.315 3.565 0.530 ;
        RECT  3.525 1.040 3.565 1.470 ;
        RECT  2.630 1.360 3.525 1.470 ;
        RECT  3.405 0.745 3.475 0.915 ;
        RECT  3.315 0.305 3.405 1.270 ;
        RECT  3.220 0.305 3.315 0.415 ;
        RECT  3.205 1.180 3.315 1.270 ;
        RECT  3.130 0.565 3.225 1.090 ;
        RECT  3.115 0.305 3.130 1.090 ;
        RECT  3.040 0.305 3.115 0.655 ;
        RECT  2.855 1.000 3.115 1.090 ;
        RECT  2.700 0.305 3.040 0.415 ;
        RECT  2.745 1.000 2.855 1.250 ;
        RECT  2.605 0.585 2.630 1.470 ;
        RECT  2.540 0.285 2.605 1.470 ;
        RECT  2.495 0.285 2.540 0.675 ;
        RECT  2.475 1.045 2.540 1.470 ;
        RECT  2.325 0.785 2.430 0.955 ;
        RECT  2.235 0.785 2.325 1.315 ;
        RECT  1.140 1.215 2.235 1.315 ;
        RECT  2.105 1.015 2.135 1.125 ;
        RECT  1.995 0.515 2.105 1.125 ;
        RECT  1.345 1.035 1.995 1.125 ;
        RECT  1.310 0.455 1.420 0.795 ;
        RECT  1.235 0.905 1.345 1.125 ;
        RECT  1.140 0.705 1.310 0.795 ;
        RECT  0.960 0.475 1.210 0.585 ;
        RECT  1.050 0.705 1.140 1.315 ;
        RECT  0.930 0.375 0.960 1.290 ;
        RECT  0.870 0.375 0.930 1.520 ;
        RECT  0.525 0.375 0.870 0.485 ;
        RECT  0.820 1.200 0.870 1.520 ;
        RECT  0.350 0.750 0.530 0.920 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.075 0.350 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.520 ;
    END
END SDFKSND4

MACRO SDFKSNQD0
    CLASS CORE ;
    FOREIGN SDFKSNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.680 0.170 1.090 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.710 2.595 0.890 ;
        RECT  2.450 0.710 2.560 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0453 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.890 ;
        RECT  1.020 0.510 1.050 0.710 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0180 ;
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.275 5.950 1.490 ;
        RECT  5.815 0.275 5.850 0.650 ;
        RECT  5.815 1.040 5.850 1.490 ;
        RECT  5.500 0.560 5.815 0.650 ;
        RECT  5.390 0.560 5.500 0.920 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.750 0.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.700 2.960 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.665 -0.165 6.000 0.165 ;
        RECT  5.555 -0.165 5.665 0.445 ;
        RECT  1.550 -0.165 5.555 0.165 ;
        RECT  1.440 -0.165 1.550 0.615 ;
        RECT  0.000 -0.165 1.440 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.625 1.635 6.000 1.965 ;
        RECT  5.515 1.415 5.625 1.965 ;
        RECT  4.480 1.635 5.515 1.965 ;
        RECT  4.370 1.385 4.480 1.965 ;
        RECT  1.465 1.635 4.370 1.965 ;
        RECT  1.355 1.475 1.465 1.965 ;
        RECT  0.475 1.635 1.355 1.965 ;
        RECT  0.305 1.385 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.750 5.750 0.920 ;
        RECT  5.615 0.750 5.705 1.305 ;
        RECT  4.970 1.195 5.615 1.305 ;
        RECT  5.170 0.975 5.285 1.085 ;
        RECT  5.060 0.275 5.170 1.085 ;
        RECT  4.925 0.275 5.060 0.365 ;
        RECT  4.880 0.480 4.970 1.305 ;
        RECT  4.715 0.255 4.925 0.365 ;
        RECT  4.860 0.480 4.880 0.675 ;
        RECT  4.770 1.105 4.790 1.315 ;
        RECT  4.680 0.505 4.770 1.315 ;
        RECT  4.190 0.275 4.715 0.365 ;
        RECT  4.360 0.505 4.680 0.620 ;
        RECT  4.480 0.730 4.590 1.295 ;
        RECT  4.015 1.190 4.480 1.295 ;
        RECT  4.250 0.505 4.360 0.940 ;
        RECT  3.975 0.255 4.190 0.365 ;
        RECT  3.905 0.465 4.015 1.295 ;
        RECT  3.835 1.190 3.905 1.295 ;
        RECT  3.475 0.795 3.765 0.925 ;
        RECT  3.615 0.275 3.735 0.485 ;
        RECT  3.615 1.070 3.725 1.525 ;
        RECT  2.010 0.275 3.615 0.365 ;
        RECT  1.970 1.435 3.615 1.525 ;
        RECT  3.375 0.475 3.475 1.290 ;
        RECT  3.160 0.720 3.285 0.890 ;
        RECT  3.070 0.465 3.160 1.290 ;
        RECT  2.820 0.465 3.070 0.575 ;
        RECT  2.810 1.180 3.070 1.290 ;
        RECT  2.355 0.465 2.730 0.575 ;
        RECT  2.355 1.180 2.720 1.290 ;
        RECT  2.245 0.465 2.355 1.290 ;
        RECT  1.985 0.725 2.095 1.105 ;
        RECT  1.900 0.275 2.010 0.615 ;
        RECT  1.350 0.725 1.985 0.815 ;
        RECT  1.860 1.215 1.970 1.525 ;
        RECT  1.680 0.950 1.885 1.060 ;
        RECT  1.590 0.950 1.680 1.375 ;
        RECT  0.930 1.285 1.590 1.375 ;
        RECT  1.240 0.305 1.350 1.175 ;
        RECT  1.115 0.305 1.240 0.415 ;
        RECT  1.025 1.065 1.240 1.175 ;
        RECT  0.895 0.305 0.930 1.375 ;
        RECT  0.840 0.305 0.895 1.515 ;
        RECT  0.525 0.305 0.840 0.415 ;
        RECT  0.785 1.285 0.840 1.515 ;
        RECT  0.350 0.870 0.570 1.005 ;
        RECT  0.260 0.480 0.350 1.290 ;
        RECT  0.185 0.480 0.260 0.570 ;
        RECT  0.185 1.200 0.260 1.290 ;
        RECT  0.075 0.300 0.185 0.570 ;
        RECT  0.075 1.200 0.185 1.515 ;
    END
END SDFKSNQD0

MACRO SDFKSNQD1
    CLASS CORE ;
    FOREIGN SDFKSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.775 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0604 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.290 2.350 0.690 ;
        RECT  2.060 0.290 2.250 0.400 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.285 6.150 1.490 ;
        RECT  6.015 0.285 6.050 0.675 ;
        RECT  6.015 1.050 6.050 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.780 0.925 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.610 0.710 2.925 0.890 ;
        RECT  2.520 0.710 2.610 1.290 ;
        RECT  2.450 1.060 2.520 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.865 -0.165 6.200 0.165 ;
        RECT  5.755 -0.165 5.865 0.685 ;
        RECT  4.285 -0.165 5.755 0.165 ;
        RECT  4.175 -0.165 4.285 0.490 ;
        RECT  1.895 -0.165 4.175 0.165 ;
        RECT  1.785 -0.165 1.895 0.400 ;
        RECT  0.000 -0.165 1.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.865 1.635 6.200 1.965 ;
        RECT  5.755 1.050 5.865 1.965 ;
        RECT  5.285 1.635 5.755 1.965 ;
        RECT  5.175 1.330 5.285 1.965 ;
        RECT  4.280 1.635 5.175 1.965 ;
        RECT  4.100 1.200 4.280 1.965 ;
        RECT  2.300 1.635 4.100 1.965 ;
        RECT  2.190 1.440 2.300 1.965 ;
        RECT  1.725 1.635 2.190 1.965 ;
        RECT  1.555 1.405 1.725 1.965 ;
        RECT  0.475 1.635 1.555 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.545 0.255 5.565 1.230 ;
        RECT  5.475 0.255 5.545 1.545 ;
        RECT  5.455 0.255 5.475 0.690 ;
        RECT  5.435 1.140 5.475 1.545 ;
        RECT  5.070 0.580 5.455 0.690 ;
        RECT  5.085 0.840 5.380 1.010 ;
        RECT  4.995 0.840 5.085 1.495 ;
        RECT  4.975 0.840 4.995 0.945 ;
        RECT  4.600 1.380 4.995 1.495 ;
        RECT  4.885 0.305 4.975 0.945 ;
        RECT  4.780 1.090 4.905 1.260 ;
        RECT  4.695 0.305 4.885 0.415 ;
        RECT  4.670 0.565 4.780 1.260 ;
        RECT  4.500 0.465 4.575 1.110 ;
        RECT  4.485 0.465 4.500 1.285 ;
        RECT  4.460 0.465 4.485 0.635 ;
        RECT  4.390 1.020 4.485 1.285 ;
        RECT  4.345 0.740 4.395 0.910 ;
        RECT  4.145 1.020 4.390 1.110 ;
        RECT  4.255 0.590 4.345 0.910 ;
        RECT  3.775 0.590 4.255 0.680 ;
        RECT  4.035 0.785 4.145 1.110 ;
        RECT  3.665 0.330 3.775 1.365 ;
        RECT  3.475 0.255 3.565 1.525 ;
        RECT  3.350 0.255 3.475 0.375 ;
        RECT  2.480 1.415 3.475 1.525 ;
        RECT  3.275 0.485 3.385 1.275 ;
        RECT  2.680 0.275 3.350 0.375 ;
        RECT  3.210 0.485 3.275 0.655 ;
        RECT  3.140 1.165 3.275 1.275 ;
        RECT  3.110 0.735 3.155 0.905 ;
        RECT  3.015 0.515 3.110 1.070 ;
        RECT  2.670 0.515 3.015 0.620 ;
        RECT  2.800 0.980 3.015 1.070 ;
        RECT  2.700 0.980 2.800 1.250 ;
        RECT  2.510 0.265 2.680 0.375 ;
        RECT  2.325 0.785 2.430 0.955 ;
        RECT  2.235 0.785 2.325 1.315 ;
        RECT  1.140 1.215 2.235 1.315 ;
        RECT  2.105 1.015 2.135 1.125 ;
        RECT  1.995 0.515 2.105 1.125 ;
        RECT  1.345 1.035 1.995 1.125 ;
        RECT  1.310 0.455 1.420 0.795 ;
        RECT  1.235 0.905 1.345 1.125 ;
        RECT  1.140 0.705 1.310 0.795 ;
        RECT  0.960 0.475 1.210 0.585 ;
        RECT  1.050 0.705 1.140 1.315 ;
        RECT  0.930 0.375 0.960 1.290 ;
        RECT  0.870 0.375 0.930 1.520 ;
        RECT  0.525 0.375 0.870 0.485 ;
        RECT  0.820 1.200 0.870 1.520 ;
        RECT  0.350 0.750 0.530 0.920 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.075 0.350 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.520 ;
    END
END SDFKSNQD1

MACRO SDFKSNQD2
    CLASS CORE ;
    FOREIGN SDFKSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.775 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0604 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.290 2.350 0.690 ;
        RECT  2.060 0.290 2.250 0.400 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.575 6.150 1.150 ;
        RECT  6.045 0.575 6.050 0.675 ;
        RECT  6.045 1.050 6.050 1.150 ;
        RECT  5.935 0.285 6.045 0.675 ;
        RECT  5.935 1.050 6.045 1.460 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.780 0.925 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.610 0.710 2.925 0.890 ;
        RECT  2.520 0.710 2.610 1.290 ;
        RECT  2.450 1.060 2.520 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.305 -0.165 6.400 0.165 ;
        RECT  6.195 -0.165 6.305 0.485 ;
        RECT  4.285 -0.165 6.195 0.165 ;
        RECT  4.175 -0.165 4.285 0.490 ;
        RECT  1.895 -0.165 4.175 0.165 ;
        RECT  1.785 -0.165 1.895 0.400 ;
        RECT  0.000 -0.165 1.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.305 1.635 6.400 1.965 ;
        RECT  6.195 1.250 6.305 1.965 ;
        RECT  5.285 1.635 6.195 1.965 ;
        RECT  5.175 1.250 5.285 1.965 ;
        RECT  4.280 1.635 5.175 1.965 ;
        RECT  4.100 1.200 4.280 1.965 ;
        RECT  2.300 1.635 4.100 1.965 ;
        RECT  2.190 1.440 2.300 1.965 ;
        RECT  1.725 1.635 2.190 1.965 ;
        RECT  1.555 1.405 1.725 1.965 ;
        RECT  0.475 1.635 1.555 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.725 0.325 5.825 1.415 ;
        RECT  5.210 0.325 5.725 0.435 ;
        RECT  5.405 1.305 5.725 1.415 ;
        RECT  5.085 0.840 5.450 1.010 ;
        RECT  5.100 0.325 5.210 0.720 ;
        RECT  4.995 0.840 5.085 1.495 ;
        RECT  4.975 0.840 4.995 0.945 ;
        RECT  4.600 1.380 4.995 1.495 ;
        RECT  4.885 0.305 4.975 0.945 ;
        RECT  4.780 1.090 4.905 1.260 ;
        RECT  4.695 0.305 4.885 0.415 ;
        RECT  4.670 0.565 4.780 1.260 ;
        RECT  4.500 0.465 4.575 1.110 ;
        RECT  4.485 0.465 4.500 1.285 ;
        RECT  4.460 0.465 4.485 0.635 ;
        RECT  4.390 1.020 4.485 1.285 ;
        RECT  4.345 0.740 4.395 0.910 ;
        RECT  4.145 1.020 4.390 1.110 ;
        RECT  4.255 0.590 4.345 0.910 ;
        RECT  3.775 0.590 4.255 0.680 ;
        RECT  4.035 0.785 4.145 1.110 ;
        RECT  3.665 0.330 3.775 1.365 ;
        RECT  3.475 0.255 3.565 1.525 ;
        RECT  3.350 0.255 3.475 0.375 ;
        RECT  2.480 1.415 3.475 1.525 ;
        RECT  3.275 0.485 3.385 1.275 ;
        RECT  2.680 0.275 3.350 0.375 ;
        RECT  3.210 0.485 3.275 0.655 ;
        RECT  3.140 1.165 3.275 1.275 ;
        RECT  3.110 0.735 3.155 0.905 ;
        RECT  3.015 0.515 3.110 1.070 ;
        RECT  2.670 0.515 3.015 0.620 ;
        RECT  2.800 0.980 3.015 1.070 ;
        RECT  2.700 0.980 2.800 1.250 ;
        RECT  2.510 0.265 2.680 0.375 ;
        RECT  2.325 0.785 2.430 0.955 ;
        RECT  2.235 0.785 2.325 1.315 ;
        RECT  1.140 1.215 2.235 1.315 ;
        RECT  2.105 1.015 2.135 1.125 ;
        RECT  1.995 0.515 2.105 1.125 ;
        RECT  1.345 1.035 1.995 1.125 ;
        RECT  1.310 0.455 1.420 0.795 ;
        RECT  1.235 0.905 1.345 1.125 ;
        RECT  1.140 0.705 1.310 0.795 ;
        RECT  0.960 0.475 1.210 0.585 ;
        RECT  1.050 0.705 1.140 1.315 ;
        RECT  0.930 0.375 0.960 1.290 ;
        RECT  0.870 0.375 0.930 1.520 ;
        RECT  0.525 0.375 0.870 0.485 ;
        RECT  0.820 1.200 0.870 1.520 ;
        RECT  0.350 0.750 0.530 0.920 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.075 0.350 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.520 ;
    END
END SDFKSNQD2

MACRO SDFKSNQD4
    CLASS CORE ;
    FOREIGN SDFKSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.170 1.100 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.510 1.775 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0604 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.290 2.350 0.690 ;
        RECT  2.060 0.290 2.250 0.400 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.355 0.295 7.465 0.675 ;
        RECT  7.355 1.020 7.465 1.470 ;
        RECT  7.250 0.525 7.355 0.675 ;
        RECT  7.250 1.020 7.355 1.190 ;
        RECT  6.950 0.525 7.250 1.190 ;
        RECT  6.945 0.525 6.950 0.675 ;
        RECT  6.835 1.020 6.950 1.490 ;
        RECT  6.835 0.295 6.945 0.675 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 0.780 0.925 ;
        RECT  0.645 0.710 0.750 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.815 0.510 2.950 0.910 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.725 -0.165 7.800 0.165 ;
        RECT  7.615 -0.165 7.725 0.695 ;
        RECT  7.235 -0.165 7.615 0.165 ;
        RECT  7.065 -0.165 7.235 0.435 ;
        RECT  4.940 -0.165 7.065 0.165 ;
        RECT  4.830 -0.165 4.940 0.685 ;
        RECT  4.325 -0.165 4.830 0.165 ;
        RECT  4.325 0.365 4.445 0.475 ;
        RECT  4.235 -0.165 4.325 0.475 ;
        RECT  1.895 -0.165 4.235 0.165 ;
        RECT  1.785 -0.165 1.895 0.400 ;
        RECT  0.000 -0.165 1.785 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.725 1.635 7.800 1.965 ;
        RECT  7.615 1.105 7.725 1.965 ;
        RECT  7.230 1.635 7.615 1.965 ;
        RECT  7.070 1.300 7.230 1.965 ;
        RECT  6.200 1.635 7.070 1.965 ;
        RECT  6.085 1.330 6.200 1.965 ;
        RECT  4.920 1.635 6.085 1.965 ;
        RECT  4.750 1.215 4.920 1.965 ;
        RECT  4.410 1.635 4.750 1.965 ;
        RECT  4.230 1.215 4.410 1.965 ;
        RECT  2.300 1.635 4.230 1.965 ;
        RECT  2.190 1.440 2.300 1.965 ;
        RECT  1.725 1.635 2.190 1.965 ;
        RECT  1.555 1.405 1.725 1.965 ;
        RECT  0.475 1.635 1.555 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.355 0.295 7.465 0.675 ;
        RECT  7.355 1.020 7.465 1.470 ;
        RECT  7.350 0.525 7.355 0.675 ;
        RECT  7.350 1.020 7.355 1.190 ;
        RECT  6.835 0.295 6.850 0.675 ;
        RECT  6.835 1.020 6.850 1.490 ;
        RECT  6.525 0.635 6.630 1.455 ;
        RECT  6.460 0.635 6.525 0.745 ;
        RECT  6.300 1.345 6.525 1.455 ;
        RECT  6.350 0.310 6.460 0.745 ;
        RECT  5.995 0.855 6.415 0.965 ;
        RECT  5.970 0.635 6.350 0.745 ;
        RECT  5.905 0.855 5.995 1.495 ;
        RECT  5.870 0.855 5.905 0.955 ;
        RECT  5.150 1.385 5.905 1.495 ;
        RECT  5.780 0.275 5.870 0.955 ;
        RECT  5.705 1.090 5.815 1.270 ;
        RECT  5.600 0.275 5.780 0.415 ;
        RECT  5.685 1.090 5.705 1.180 ;
        RECT  5.575 0.560 5.685 1.180 ;
        RECT  5.190 0.275 5.600 0.365 ;
        RECT  5.410 0.455 5.475 0.625 ;
        RECT  5.320 0.455 5.410 1.270 ;
        RECT  5.300 0.790 5.320 1.270 ;
        RECT  4.705 0.790 5.300 0.880 ;
        RECT  5.080 0.275 5.190 0.465 ;
        RECT  5.040 1.045 5.150 1.495 ;
        RECT  4.630 0.465 4.705 1.110 ;
        RECT  4.615 0.465 4.630 1.285 ;
        RECT  4.570 0.465 4.615 0.635 ;
        RECT  4.520 1.020 4.615 1.285 ;
        RECT  4.445 0.740 4.525 0.910 ;
        RECT  4.265 1.020 4.520 1.110 ;
        RECT  4.355 0.575 4.445 0.910 ;
        RECT  3.885 0.575 4.355 0.665 ;
        RECT  4.165 0.775 4.265 1.110 ;
        RECT  3.775 0.325 3.885 1.365 ;
        RECT  3.565 0.315 3.655 1.470 ;
        RECT  3.515 0.315 3.565 0.530 ;
        RECT  3.525 1.040 3.565 1.470 ;
        RECT  2.630 1.360 3.525 1.470 ;
        RECT  3.405 0.745 3.475 0.915 ;
        RECT  3.315 0.305 3.405 1.270 ;
        RECT  3.220 0.305 3.315 0.415 ;
        RECT  3.205 1.180 3.315 1.270 ;
        RECT  3.130 0.565 3.225 1.090 ;
        RECT  3.115 0.305 3.130 1.090 ;
        RECT  3.040 0.305 3.115 0.655 ;
        RECT  2.855 1.000 3.115 1.090 ;
        RECT  2.700 0.305 3.040 0.415 ;
        RECT  2.745 1.000 2.855 1.250 ;
        RECT  2.605 0.585 2.630 1.470 ;
        RECT  2.540 0.285 2.605 1.470 ;
        RECT  2.495 0.285 2.540 0.675 ;
        RECT  2.475 1.045 2.540 1.470 ;
        RECT  2.325 0.785 2.430 0.955 ;
        RECT  2.235 0.785 2.325 1.315 ;
        RECT  1.140 1.215 2.235 1.315 ;
        RECT  2.105 1.015 2.135 1.125 ;
        RECT  1.995 0.515 2.105 1.125 ;
        RECT  1.345 1.035 1.995 1.125 ;
        RECT  1.310 0.455 1.420 0.795 ;
        RECT  1.235 0.905 1.345 1.125 ;
        RECT  1.140 0.705 1.310 0.795 ;
        RECT  0.960 0.475 1.210 0.585 ;
        RECT  1.050 0.705 1.140 1.315 ;
        RECT  0.930 0.375 0.960 1.290 ;
        RECT  0.870 0.375 0.930 1.520 ;
        RECT  0.525 0.375 0.870 0.485 ;
        RECT  0.820 1.200 0.870 1.520 ;
        RECT  0.350 0.750 0.530 0.920 ;
        RECT  0.260 0.500 0.350 1.300 ;
        RECT  0.185 0.500 0.260 0.590 ;
        RECT  0.185 1.210 0.260 1.300 ;
        RECT  0.075 0.350 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.520 ;
    END
END SDFKSNQD4

MACRO SDFNCND0
    CLASS CORE ;
    FOREIGN SDFNCND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.485 6.150 1.490 ;
        RECT  6.020 0.485 6.050 0.675 ;
        RECT  6.010 1.280 6.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.505 5.750 1.440 ;
        RECT  5.475 0.505 5.650 0.615 ;
        RECT  5.460 1.330 5.650 1.440 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.880 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0667 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.005 0.910 5.150 1.090 ;
        RECT  4.850 0.845 5.005 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.825 -0.165 6.200 0.165 ;
        RECT  4.655 -0.165 4.825 0.355 ;
        RECT  3.520 -0.165 4.655 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.635 6.200 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.930 0.750 5.960 0.920 ;
        RECT  5.840 0.275 5.930 0.920 ;
        RECT  5.080 0.275 5.840 0.365 ;
        RECT  5.370 0.735 5.560 0.845 ;
        RECT  5.350 1.015 5.540 1.125 ;
        RECT  5.270 0.455 5.370 0.845 ;
        RECT  5.260 1.015 5.350 1.525 ;
        RECT  5.250 0.455 5.270 0.715 ;
        RECT  4.315 1.435 5.260 1.525 ;
        RECT  4.755 0.625 5.250 0.715 ;
        RECT  4.755 1.225 5.150 1.335 ;
        RECT  4.990 0.275 5.080 0.535 ;
        RECT  4.575 0.445 4.990 0.535 ;
        RECT  4.665 0.625 4.755 1.335 ;
        RECT  4.485 0.445 4.575 1.335 ;
        RECT  4.410 0.445 4.485 0.640 ;
        RECT  4.405 1.225 4.485 1.335 ;
        RECT  4.320 0.750 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  4.230 0.315 4.285 0.840 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.820 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.460 0.275 2.570 0.445 ;
        RECT  0.865 0.305 2.460 0.405 ;
        RECT  2.305 1.295 2.405 1.525 ;
        RECT  2.230 0.495 2.350 1.135 ;
        RECT  0.945 1.295 2.305 1.385 ;
        RECT  2.110 0.495 2.230 0.605 ;
        RECT  2.065 1.025 2.230 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.500 1.960 1.195 ;
        RECT  1.615 0.500 1.860 0.610 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.260 0.500 1.360 0.845 ;
        RECT  0.850 0.500 1.260 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.500 0.850 0.915 ;
        RECT  0.355 0.500 0.740 0.590 ;
        RECT  0.265 0.500 0.355 1.290 ;
        RECT  0.185 0.500 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNCND0

MACRO SDFNCND1
    CLASS CORE ;
    FOREIGN SDFNCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.025 ;
        RECT  0.445 0.680 0.555 1.320 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.680 0.355 1.120 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1480 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.275 6.150 1.490 ;
        RECT  6.020 0.275 6.050 0.675 ;
        RECT  6.010 1.080 6.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.505 5.750 1.440 ;
        RECT  5.475 0.505 5.650 0.615 ;
        RECT  5.460 1.330 5.650 1.440 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.785 1.610 0.975 ;
        RECT  1.445 0.495 1.555 0.975 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0667 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.005 0.910 5.150 1.090 ;
        RECT  4.850 0.845 5.005 1.090 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.825 -0.165 6.200 0.165 ;
        RECT  4.655 -0.165 4.825 0.355 ;
        RECT  3.520 -0.165 4.655 0.165 ;
        RECT  3.410 -0.165 3.520 0.415 ;
        RECT  0.520 -0.165 3.410 0.165 ;
        RECT  0.310 -0.165 0.520 0.370 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.635 6.200 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.610 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.610 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.520 1.635 1.570 1.965 ;
        RECT  0.310 1.430 0.520 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.930 0.750 5.960 0.920 ;
        RECT  5.840 0.275 5.930 0.920 ;
        RECT  5.080 0.275 5.840 0.365 ;
        RECT  5.370 0.735 5.560 0.845 ;
        RECT  5.350 1.015 5.540 1.125 ;
        RECT  5.270 0.455 5.370 0.845 ;
        RECT  5.260 1.015 5.350 1.525 ;
        RECT  5.250 0.455 5.270 0.715 ;
        RECT  4.315 1.435 5.260 1.525 ;
        RECT  4.755 0.625 5.250 0.715 ;
        RECT  4.755 1.225 5.150 1.335 ;
        RECT  4.990 0.275 5.080 0.535 ;
        RECT  4.575 0.445 4.990 0.535 ;
        RECT  4.665 0.625 4.755 1.335 ;
        RECT  4.485 0.445 4.575 1.335 ;
        RECT  4.410 0.445 4.485 0.640 ;
        RECT  4.405 1.225 4.485 1.335 ;
        RECT  4.320 0.750 4.395 1.120 ;
        RECT  4.285 0.315 4.320 1.120 ;
        RECT  4.225 1.225 4.315 1.525 ;
        RECT  4.230 0.315 4.285 0.840 ;
        RECT  3.700 0.315 4.230 0.415 ;
        RECT  4.140 1.225 4.225 1.335 ;
        RECT  4.050 0.505 4.140 1.335 ;
        RECT  3.945 1.435 4.135 1.545 ;
        RECT  4.030 0.505 4.050 0.705 ;
        RECT  3.900 1.125 3.960 1.320 ;
        RECT  2.890 1.435 3.945 1.525 ;
        RECT  3.850 0.505 3.900 1.320 ;
        RECT  3.790 0.505 3.850 1.225 ;
        RECT  3.485 1.125 3.790 1.225 ;
        RECT  3.610 0.315 3.700 0.595 ;
        RECT  3.590 0.685 3.700 0.940 ;
        RECT  3.230 0.505 3.610 0.595 ;
        RECT  2.875 0.685 3.590 0.785 ;
        RECT  3.385 0.910 3.485 1.225 ;
        RECT  2.970 0.910 3.385 1.030 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.820 0.275 3.130 0.365 ;
        RECT  2.700 1.435 2.890 1.545 ;
        RECT  2.860 0.455 2.875 0.785 ;
        RECT  2.765 0.455 2.860 1.155 ;
        RECT  2.565 1.045 2.765 1.155 ;
        RECT  2.460 0.275 2.570 0.445 ;
        RECT  0.865 0.315 2.460 0.405 ;
        RECT  2.305 1.295 2.405 1.525 ;
        RECT  2.230 0.495 2.350 1.135 ;
        RECT  1.460 1.295 2.305 1.385 ;
        RECT  2.110 0.495 2.230 0.605 ;
        RECT  2.065 1.025 2.230 1.135 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.515 1.960 1.195 ;
        RECT  1.675 0.515 1.860 0.685 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.500 ;
        RECT  0.940 1.410 1.360 1.500 ;
        RECT  1.140 0.500 1.325 0.590 ;
        RECT  1.140 1.210 1.250 1.310 ;
        RECT  1.050 0.500 1.140 1.310 ;
        RECT  0.835 1.135 0.940 1.500 ;
        RECT  0.750 0.595 0.840 0.925 ;
        RECT  0.730 0.460 0.750 0.925 ;
        RECT  0.660 0.460 0.730 0.705 ;
        RECT  0.185 0.460 0.660 0.570 ;
        RECT  0.150 0.400 0.185 0.570 ;
        RECT  0.150 1.230 0.185 1.460 ;
        RECT  0.060 0.400 0.150 1.460 ;
    END
END SDFNCND1

MACRO SDFNCND2
    CLASS CORE ;
    FOREIGN SDFNCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.025 ;
        RECT  0.445 0.680 0.555 1.320 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.680 0.355 1.120 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.685 0.510 6.750 1.310 ;
        RECT  6.645 0.285 6.685 1.490 ;
        RECT  6.565 0.285 6.645 0.660 ;
        RECT  6.560 1.080 6.645 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.080 0.485 6.175 1.490 ;
        RECT  6.045 0.485 6.080 0.660 ;
        RECT  6.045 1.025 6.080 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.785 1.610 0.975 ;
        RECT  1.445 0.495 1.555 0.975 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0877 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.640 0.710 5.755 1.135 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.955 -0.165 7.000 0.165 ;
        RECT  4.785 -0.165 4.955 0.355 ;
        RECT  3.530 -0.165 4.785 0.165 ;
        RECT  3.420 -0.165 3.530 0.405 ;
        RECT  0.520 -0.165 3.420 0.165 ;
        RECT  0.310 -0.165 0.520 0.370 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.580 1.635 7.000 1.965 ;
        RECT  3.580 1.215 3.750 1.305 ;
        RECT  3.470 1.215 3.580 1.965 ;
        RECT  3.175 1.635 3.470 1.965 ;
        RECT  3.175 1.125 3.285 1.235 ;
        RECT  3.085 1.125 3.175 1.965 ;
        RECT  1.760 1.635 3.085 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.520 1.635 1.570 1.965 ;
        RECT  0.310 1.430 0.520 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.420 0.750 6.510 0.920 ;
        RECT  6.330 0.280 6.420 0.920 ;
        RECT  5.175 0.280 6.330 0.370 ;
        RECT  5.935 0.750 5.990 0.920 ;
        RECT  5.845 0.495 5.935 1.420 ;
        RECT  5.375 0.495 5.845 0.600 ;
        RECT  5.485 1.285 5.845 1.420 ;
        RECT  5.355 0.950 5.460 1.060 ;
        RECT  5.285 0.495 5.375 0.810 ;
        RECT  5.265 0.950 5.355 1.525 ;
        RECT  4.880 0.720 5.285 0.810 ;
        RECT  4.325 1.435 5.265 1.525 ;
        RECT  5.085 0.280 5.175 0.545 ;
        RECT  4.880 1.215 5.140 1.325 ;
        RECT  4.655 0.455 5.085 0.545 ;
        RECT  4.770 0.720 4.880 1.325 ;
        RECT  4.565 0.455 4.655 1.345 ;
        RECT  4.480 0.455 4.565 0.695 ;
        RECT  4.435 1.245 4.565 1.345 ;
        RECT  4.390 0.945 4.475 1.115 ;
        RECT  4.300 0.325 4.390 1.115 ;
        RECT  4.230 1.245 4.325 1.525 ;
        RECT  3.730 0.325 4.300 0.415 ;
        RECT  4.200 1.245 4.230 1.355 ;
        RECT  4.090 0.505 4.200 1.355 ;
        RECT  3.870 0.505 3.970 1.335 ;
        RECT  3.840 0.505 3.870 0.675 ;
        RECT  3.465 1.035 3.870 1.125 ;
        RECT  3.630 0.685 3.740 0.905 ;
        RECT  3.640 0.325 3.730 0.585 ;
        RECT  3.230 0.495 3.640 0.585 ;
        RECT  2.820 0.685 3.630 0.785 ;
        RECT  3.375 0.895 3.465 1.125 ;
        RECT  2.970 0.895 3.375 1.005 ;
        RECT  3.130 0.275 3.230 0.585 ;
        RECT  2.765 0.275 3.130 0.365 ;
        RECT  2.710 0.465 2.820 1.165 ;
        RECT  2.695 1.040 2.710 1.165 ;
        RECT  2.585 1.040 2.695 1.505 ;
        RECT  2.450 0.315 2.560 0.645 ;
        RECT  0.865 0.315 2.450 0.405 ;
        RECT  2.285 1.295 2.405 1.515 ;
        RECT  2.240 0.495 2.340 1.155 ;
        RECT  1.460 1.295 2.285 1.385 ;
        RECT  2.110 0.495 2.240 0.585 ;
        RECT  2.045 1.045 2.240 1.155 ;
        RECT  1.935 0.760 2.085 0.930 ;
        RECT  1.825 0.515 1.935 1.195 ;
        RECT  1.675 0.515 1.825 0.685 ;
        RECT  1.555 1.085 1.825 1.195 ;
        RECT  1.360 1.295 1.460 1.500 ;
        RECT  0.940 1.410 1.360 1.500 ;
        RECT  1.140 0.500 1.325 0.590 ;
        RECT  1.140 1.210 1.250 1.310 ;
        RECT  1.050 0.500 1.140 1.310 ;
        RECT  0.835 1.135 0.940 1.500 ;
        RECT  0.750 0.595 0.840 0.925 ;
        RECT  0.730 0.460 0.750 0.925 ;
        RECT  0.660 0.460 0.730 0.705 ;
        RECT  0.185 0.460 0.660 0.570 ;
        RECT  0.150 0.400 0.185 0.570 ;
        RECT  0.150 1.230 0.185 1.460 ;
        RECT  0.060 0.400 0.150 1.460 ;
    END
END SDFNCND2

MACRO SDFNCND4
    CLASS CORE ;
    FOREIGN SDFNCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.025 ;
        RECT  0.445 0.680 0.555 1.320 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.680 0.355 1.120 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 0.325 8.150 0.635 ;
        RECT  8.050 1.100 8.150 1.410 ;
        RECT  7.750 0.325 8.050 1.410 ;
        RECT  7.435 0.325 7.750 0.635 ;
        RECT  7.435 1.100 7.750 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 1.100 7.150 1.410 ;
        RECT  7.050 0.510 7.105 0.690 ;
        RECT  6.750 0.510 7.050 1.410 ;
        RECT  6.435 0.510 6.750 0.695 ;
        RECT  6.435 1.100 6.750 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.700 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.775 1.610 0.975 ;
        RECT  1.445 0.495 1.555 0.975 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0876 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.550 0.965 5.685 1.135 ;
        RECT  5.450 0.710 5.550 1.135 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.915 -0.165 8.400 0.165 ;
        RECT  4.745 -0.165 4.915 0.355 ;
        RECT  3.530 -0.165 4.745 0.165 ;
        RECT  3.420 -0.165 3.530 0.405 ;
        RECT  0.520 -0.165 3.420 0.165 ;
        RECT  0.310 -0.165 0.520 0.370 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 1.635 8.400 1.965 ;
        RECT  3.610 1.175 3.720 1.965 ;
        RECT  3.175 1.635 3.610 1.965 ;
        RECT  3.175 1.130 3.285 1.240 ;
        RECT  3.085 1.130 3.175 1.965 ;
        RECT  0.520 1.635 3.085 1.965 ;
        RECT  0.310 1.430 0.520 1.965 ;
        RECT  0.000 1.635 0.310 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.435 0.325 7.650 0.635 ;
        RECT  7.435 1.100 7.650 1.410 ;
        RECT  6.435 0.510 6.650 0.695 ;
        RECT  6.435 1.100 6.650 1.410 ;
        RECT  7.320 0.775 7.500 0.895 ;
        RECT  7.230 0.280 7.320 0.895 ;
        RECT  6.305 0.280 7.230 0.370 ;
        RECT  6.215 0.280 6.305 1.170 ;
        RECT  6.075 0.280 6.215 0.370 ;
        RECT  6.075 1.080 6.215 1.170 ;
        RECT  5.975 0.280 6.075 0.650 ;
        RECT  5.975 1.080 6.075 1.460 ;
        RECT  5.880 0.760 6.050 0.930 ;
        RECT  5.120 0.280 5.975 0.370 ;
        RECT  5.790 0.495 5.880 1.410 ;
        RECT  5.320 0.495 5.790 0.600 ;
        RECT  5.460 1.300 5.790 1.410 ;
        RECT  5.230 0.920 5.340 1.525 ;
        RECT  5.230 0.495 5.320 0.810 ;
        RECT  4.815 0.720 5.230 0.810 ;
        RECT  4.325 1.435 5.230 1.525 ;
        RECT  4.815 1.215 5.140 1.325 ;
        RECT  5.030 0.280 5.120 0.545 ;
        RECT  4.625 0.455 5.030 0.545 ;
        RECT  4.715 0.720 4.815 1.325 ;
        RECT  4.535 0.455 4.625 1.325 ;
        RECT  4.440 0.455 4.535 0.635 ;
        RECT  4.435 1.215 4.535 1.325 ;
        RECT  4.350 0.945 4.445 1.115 ;
        RECT  4.260 0.325 4.350 1.115 ;
        RECT  4.215 1.215 4.325 1.525 ;
        RECT  3.730 0.325 4.260 0.415 ;
        RECT  4.170 1.215 4.215 1.325 ;
        RECT  4.060 0.505 4.170 1.325 ;
        RECT  3.870 0.505 3.970 1.335 ;
        RECT  3.820 0.505 3.870 0.675 ;
        RECT  3.465 0.995 3.870 1.085 ;
        RECT  3.640 0.325 3.730 0.585 ;
        RECT  3.635 0.685 3.730 0.885 ;
        RECT  3.230 0.495 3.640 0.585 ;
        RECT  2.820 0.685 3.635 0.785 ;
        RECT  3.375 0.895 3.465 1.085 ;
        RECT  2.970 0.895 3.375 1.005 ;
        RECT  3.130 0.275 3.230 0.585 ;
        RECT  2.765 0.275 3.130 0.365 ;
        RECT  2.710 0.465 2.820 1.165 ;
        RECT  2.695 1.040 2.710 1.165 ;
        RECT  2.585 1.040 2.695 1.505 ;
        RECT  2.450 0.315 2.560 0.645 ;
        RECT  0.940 1.410 2.485 1.500 ;
        RECT  0.865 0.315 2.450 0.405 ;
        RECT  2.240 0.495 2.340 1.155 ;
        RECT  2.100 0.495 2.240 0.585 ;
        RECT  2.045 1.045 2.240 1.155 ;
        RECT  1.910 0.760 2.085 0.930 ;
        RECT  1.800 0.515 1.910 1.295 ;
        RECT  1.675 0.515 1.800 0.685 ;
        RECT  1.555 1.150 1.800 1.295 ;
        RECT  1.140 0.500 1.325 0.590 ;
        RECT  1.140 1.210 1.250 1.310 ;
        RECT  1.050 0.500 1.140 1.310 ;
        RECT  0.835 1.135 0.940 1.500 ;
        RECT  0.750 0.595 0.840 0.930 ;
        RECT  0.730 0.460 0.750 0.930 ;
        RECT  0.660 0.460 0.730 0.705 ;
        RECT  0.185 0.460 0.660 0.570 ;
        RECT  0.150 0.400 0.185 0.570 ;
        RECT  0.150 1.230 0.185 1.460 ;
        RECT  0.060 0.400 0.150 1.460 ;
    END
END SDFNCND4

MACRO SDFNCSND0
    CLASS CORE ;
    FOREIGN SDFNCSND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0583 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.710 6.150 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.825 0.475 6.950 1.330 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.530 6.550 1.295 ;
        RECT  6.260 0.530 6.450 0.640 ;
        RECT  6.260 1.185 6.450 1.295 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0355 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  1.000 0.710 1.050 0.920 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 7.000 0.165 ;
        RECT  3.420 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.420 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.620 1.635 7.000 1.965 ;
        RECT  5.450 1.400 5.620 1.965 ;
        RECT  5.050 1.635 5.450 1.965 ;
        RECT  4.880 1.405 5.050 1.965 ;
        RECT  2.590 1.635 4.880 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.590 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.590 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.645 0.275 6.735 1.515 ;
        RECT  6.105 0.275 6.645 0.375 ;
        RECT  5.910 1.405 6.645 1.515 ;
        RECT  6.240 0.750 6.350 1.090 ;
        RECT  5.760 1.000 6.240 1.090 ;
        RECT  5.995 0.275 6.105 0.465 ;
        RECT  4.860 0.275 5.995 0.365 ;
        RECT  5.800 1.180 5.910 1.515 ;
        RECT  5.710 0.455 5.760 1.090 ;
        RECT  5.660 0.455 5.710 1.290 ;
        RECT  4.950 0.455 5.660 0.565 ;
        RECT  5.620 1.005 5.660 1.290 ;
        RECT  5.165 1.180 5.620 1.290 ;
        RECT  5.440 0.710 5.530 1.090 ;
        RECT  5.045 1.000 5.440 1.090 ;
        RECT  4.955 1.000 5.045 1.305 ;
        RECT  4.510 1.215 4.955 1.305 ;
        RECT  4.770 0.275 4.860 1.125 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.410 0.980 4.510 1.305 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.700 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.465 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.820 0.685 3.605 0.785 ;
        RECT  3.375 0.895 3.465 1.295 ;
        RECT  2.970 0.895 3.375 1.005 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.765 0.275 3.130 0.375 ;
        RECT  2.710 0.465 2.820 1.165 ;
        RECT  2.540 1.065 2.710 1.165 ;
        RECT  2.450 0.305 2.560 0.645 ;
        RECT  0.865 0.305 2.450 0.405 ;
        RECT  2.295 1.295 2.405 1.525 ;
        RECT  2.240 0.510 2.340 1.135 ;
        RECT  0.945 1.295 2.295 1.385 ;
        RECT  2.110 0.510 2.240 0.620 ;
        RECT  2.065 1.025 2.240 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.500 1.960 1.195 ;
        RECT  1.615 0.500 1.860 0.610 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.255 0.495 1.360 0.845 ;
        RECT  0.850 0.495 1.255 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.495 0.850 0.915 ;
        RECT  0.355 0.495 0.740 0.590 ;
        RECT  0.265 0.495 0.355 1.290 ;
        RECT  0.185 0.495 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.460 ;
    END
END SDFNCSND0

MACRO SDFNCSND1
    CLASS CORE ;
    FOREIGN SDFNCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0646 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.710 6.150 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.825 0.285 6.950 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.525 6.550 1.295 ;
        RECT  6.260 0.525 6.450 0.635 ;
        RECT  6.260 1.185 6.450 1.295 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 7.000 0.165 ;
        RECT  3.420 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.420 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.620 1.635 7.000 1.965 ;
        RECT  5.450 1.400 5.620 1.965 ;
        RECT  5.050 1.635 5.450 1.965 ;
        RECT  4.880 1.405 5.050 1.965 ;
        RECT  2.590 1.635 4.880 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.590 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.590 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.645 0.275 6.735 1.515 ;
        RECT  6.105 0.275 6.645 0.375 ;
        RECT  5.910 1.405 6.645 1.515 ;
        RECT  6.240 0.750 6.350 1.095 ;
        RECT  5.760 1.005 6.240 1.095 ;
        RECT  5.995 0.275 6.105 0.500 ;
        RECT  4.860 0.275 5.995 0.365 ;
        RECT  5.800 1.185 5.910 1.515 ;
        RECT  5.710 0.455 5.760 1.095 ;
        RECT  5.660 0.455 5.710 1.290 ;
        RECT  4.950 0.455 5.660 0.565 ;
        RECT  5.620 1.005 5.660 1.290 ;
        RECT  5.165 1.180 5.620 1.290 ;
        RECT  5.440 0.710 5.530 1.090 ;
        RECT  5.045 1.000 5.440 1.090 ;
        RECT  4.955 1.000 5.045 1.305 ;
        RECT  4.510 1.215 4.955 1.305 ;
        RECT  4.770 0.275 4.860 1.125 ;
        RECT  4.600 0.440 4.770 0.610 ;
        RECT  4.665 1.015 4.770 1.125 ;
        RECT  4.575 0.725 4.680 0.905 ;
        RECT  4.510 0.725 4.575 0.815 ;
        RECT  4.420 0.315 4.510 0.815 ;
        RECT  4.410 0.980 4.510 1.305 ;
        RECT  4.285 1.395 4.465 1.525 ;
        RECT  3.730 0.315 4.420 0.415 ;
        RECT  4.330 0.980 4.410 1.070 ;
        RECT  4.220 0.505 4.330 1.070 ;
        RECT  3.940 1.185 4.300 1.295 ;
        RECT  2.700 1.435 4.285 1.525 ;
        RECT  3.940 0.530 4.130 0.640 ;
        RECT  3.850 0.530 3.940 1.295 ;
        RECT  3.465 1.185 3.850 1.295 ;
        RECT  3.640 0.315 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.820 0.685 3.605 0.785 ;
        RECT  3.375 0.895 3.465 1.295 ;
        RECT  2.970 0.895 3.375 1.005 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.765 0.275 3.130 0.375 ;
        RECT  2.710 0.465 2.820 1.165 ;
        RECT  2.540 1.065 2.710 1.165 ;
        RECT  2.450 0.305 2.560 0.645 ;
        RECT  0.865 0.305 2.450 0.405 ;
        RECT  2.295 1.295 2.405 1.525 ;
        RECT  2.240 0.510 2.340 1.135 ;
        RECT  1.460 1.295 2.295 1.385 ;
        RECT  2.110 0.510 2.240 0.620 ;
        RECT  2.065 1.025 2.240 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNCSND1

MACRO SDFNCSND2
    CLASS CORE ;
    FOREIGN SDFNCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0646 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.970 0.710 6.010 0.890 ;
        RECT  5.850 0.510 5.970 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.285 7.150 1.490 ;
        RECT  6.965 0.285 7.050 0.675 ;
        RECT  6.965 1.060 7.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.550 0.465 6.575 0.675 ;
        RECT  6.550 1.030 6.575 1.240 ;
        RECT  6.450 0.465 6.550 1.240 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0630 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.350 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 -0.165 7.400 0.165 ;
        RECT  3.420 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.420 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.265 1.635 7.400 1.965 ;
        RECT  6.095 1.510 6.265 1.965 ;
        RECT  5.620 1.635 6.095 1.965 ;
        RECT  5.450 1.400 5.620 1.965 ;
        RECT  5.050 1.635 5.450 1.965 ;
        RECT  4.880 1.405 5.050 1.965 ;
        RECT  2.590 1.635 4.880 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.590 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.590 1.965 ;
        RECT  1.760 1.635 2.500 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.800 0.780 6.960 0.890 ;
        RECT  6.710 0.275 6.800 1.420 ;
        RECT  6.135 0.275 6.710 0.375 ;
        RECT  5.910 1.330 6.710 1.420 ;
        RECT  6.220 0.750 6.330 1.095 ;
        RECT  5.760 1.005 6.220 1.095 ;
        RECT  5.920 0.275 6.135 0.420 ;
        RECT  4.860 0.275 5.920 0.365 ;
        RECT  5.800 1.185 5.910 1.420 ;
        RECT  5.710 0.455 5.760 1.095 ;
        RECT  5.660 0.455 5.710 1.290 ;
        RECT  4.950 0.455 5.660 0.565 ;
        RECT  5.620 1.005 5.660 1.290 ;
        RECT  5.165 1.180 5.620 1.290 ;
        RECT  5.440 0.710 5.530 1.090 ;
        RECT  5.045 1.000 5.440 1.090 ;
        RECT  4.955 1.000 5.045 1.295 ;
        RECT  4.520 1.205 4.955 1.295 ;
        RECT  4.765 0.275 4.860 1.115 ;
        RECT  4.600 0.440 4.765 0.610 ;
        RECT  4.650 1.015 4.765 1.115 ;
        RECT  4.565 0.745 4.675 0.915 ;
        RECT  4.510 0.745 4.565 0.835 ;
        RECT  4.410 1.005 4.520 1.295 ;
        RECT  4.420 0.325 4.510 0.835 ;
        RECT  4.275 1.385 4.465 1.525 ;
        RECT  3.730 0.325 4.420 0.415 ;
        RECT  4.330 1.005 4.410 1.095 ;
        RECT  4.220 0.505 4.330 1.095 ;
        RECT  3.940 1.185 4.300 1.275 ;
        RECT  2.700 1.435 4.275 1.525 ;
        RECT  3.940 0.540 4.105 0.650 ;
        RECT  3.850 0.540 3.940 1.275 ;
        RECT  3.465 1.165 3.850 1.275 ;
        RECT  3.640 0.325 3.730 0.595 ;
        RECT  3.555 0.685 3.655 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.820 0.685 3.555 0.785 ;
        RECT  3.375 0.895 3.465 1.275 ;
        RECT  2.970 0.895 3.375 1.005 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.765 0.275 3.130 0.365 ;
        RECT  2.710 0.465 2.820 1.165 ;
        RECT  2.540 1.065 2.710 1.165 ;
        RECT  2.450 0.305 2.560 0.645 ;
        RECT  0.865 0.305 2.450 0.405 ;
        RECT  2.295 1.295 2.405 1.525 ;
        RECT  2.240 0.510 2.340 1.135 ;
        RECT  1.460 1.295 2.295 1.385 ;
        RECT  2.110 0.510 2.240 0.620 ;
        RECT  2.065 1.025 2.240 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNCSND2

MACRO SDFNCSND4
    CLASS CORE ;
    FOREIGN SDFNCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0811 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.710 6.550 0.890 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.450 0.315 8.550 0.645 ;
        RECT  8.450 1.090 8.550 1.420 ;
        RECT  8.150 0.315 8.450 1.420 ;
        RECT  7.835 0.315 8.150 0.645 ;
        RECT  7.835 1.090 8.150 1.420 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.505 7.505 0.675 ;
        RECT  7.250 1.070 7.505 1.240 ;
        RECT  6.950 0.505 7.250 1.240 ;
        RECT  6.835 0.505 6.950 0.675 ;
        RECT  6.835 1.070 6.950 1.240 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0895 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.710 5.550 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.040 -0.165 8.800 0.165 ;
        RECT  4.950 -0.165 5.040 0.410 ;
        RECT  3.530 -0.165 4.950 0.165 ;
        RECT  3.420 -0.165 3.530 0.415 ;
        RECT  0.520 -0.165 3.420 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 1.635 8.800 1.965 ;
        RECT  6.495 1.510 6.665 1.965 ;
        RECT  5.040 1.635 6.495 1.965 ;
        RECT  4.870 1.405 5.040 1.965 ;
        RECT  2.590 1.635 4.870 1.965 ;
        RECT  3.090 1.125 3.285 1.235 ;
        RECT  3.000 1.125 3.090 1.345 ;
        RECT  2.590 1.255 3.000 1.345 ;
        RECT  2.500 1.255 2.590 1.965 ;
        RECT  0.470 1.635 2.500 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.835 0.315 8.050 0.645 ;
        RECT  7.835 1.090 8.050 1.420 ;
        RECT  7.350 0.505 7.505 0.675 ;
        RECT  7.350 1.070 7.505 1.240 ;
        RECT  6.835 0.505 6.850 0.675 ;
        RECT  6.835 1.070 6.850 1.240 ;
        RECT  7.700 0.780 7.920 0.890 ;
        RECT  7.610 0.275 7.700 1.420 ;
        RECT  6.495 0.275 7.610 0.375 ;
        RECT  6.330 1.330 7.610 1.420 ;
        RECT  6.640 0.730 6.745 1.095 ;
        RECT  6.150 1.005 6.640 1.095 ;
        RECT  6.385 0.275 6.495 0.585 ;
        RECT  5.220 0.275 6.385 0.365 ;
        RECT  6.220 1.185 6.330 1.420 ;
        RECT  6.130 0.485 6.150 1.095 ;
        RECT  6.040 0.485 6.130 1.270 ;
        RECT  5.425 0.485 6.040 0.595 ;
        RECT  5.155 1.160 6.040 1.270 ;
        RECT  5.800 0.710 5.910 1.070 ;
        RECT  5.160 0.980 5.800 1.070 ;
        RECT  5.130 0.275 5.220 0.610 ;
        RECT  5.050 0.710 5.160 1.070 ;
        RECT  4.860 0.520 5.130 0.610 ;
        RECT  5.045 0.980 5.050 1.070 ;
        RECT  4.955 0.980 5.045 1.295 ;
        RECT  4.520 1.205 4.955 1.295 ;
        RECT  4.765 0.435 4.860 1.115 ;
        RECT  4.600 0.435 4.765 0.610 ;
        RECT  4.650 1.015 4.765 1.115 ;
        RECT  4.565 0.745 4.675 0.915 ;
        RECT  4.510 0.745 4.565 0.835 ;
        RECT  4.410 1.005 4.520 1.295 ;
        RECT  4.420 0.325 4.510 0.835 ;
        RECT  4.275 1.385 4.465 1.525 ;
        RECT  3.730 0.325 4.420 0.415 ;
        RECT  4.330 1.005 4.410 1.095 ;
        RECT  4.220 0.505 4.330 1.095 ;
        RECT  3.940 1.185 4.300 1.275 ;
        RECT  2.700 1.435 4.275 1.525 ;
        RECT  3.940 0.540 4.120 0.650 ;
        RECT  3.850 0.540 3.940 1.275 ;
        RECT  3.465 1.165 3.850 1.275 ;
        RECT  3.640 0.325 3.730 0.595 ;
        RECT  3.605 0.685 3.715 1.025 ;
        RECT  3.230 0.505 3.640 0.595 ;
        RECT  2.820 0.685 3.605 0.785 ;
        RECT  3.375 0.895 3.465 1.275 ;
        RECT  2.970 0.895 3.375 1.005 ;
        RECT  3.130 0.275 3.230 0.595 ;
        RECT  2.765 0.275 3.130 0.365 ;
        RECT  2.710 0.465 2.820 1.165 ;
        RECT  2.560 1.055 2.710 1.165 ;
        RECT  2.450 0.305 2.560 0.645 ;
        RECT  0.865 0.305 2.450 0.405 ;
        RECT  2.305 1.325 2.405 1.525 ;
        RECT  2.235 0.510 2.345 1.165 ;
        RECT  0.945 1.435 2.305 1.525 ;
        RECT  2.110 0.510 2.235 0.620 ;
        RECT  2.065 1.055 2.235 1.165 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.325 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.215 1.860 1.325 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNCSND4

MACRO SDFND0
    CLASS CORE ;
    FOREIGN SDFND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.485 5.350 1.290 ;
        RECT  5.215 0.485 5.250 0.665 ;
        RECT  5.215 1.035 5.250 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.455 4.575 0.645 ;
        RECT  4.550 1.045 4.565 1.290 ;
        RECT  4.450 0.455 4.550 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.880 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.400 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 1.635 5.400 1.965 ;
        RECT  5.000 1.455 5.110 1.965 ;
        RECT  3.120 1.635 5.000 1.965 ;
        RECT  3.010 1.385 3.120 1.965 ;
        RECT  1.760 1.635 3.010 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.750 5.160 0.920 ;
        RECT  4.985 0.275 5.075 0.920 ;
        RECT  4.340 0.275 4.985 0.365 ;
        RECT  4.710 0.455 4.825 1.245 ;
        RECT  3.685 1.395 4.745 1.505 ;
        RECT  4.650 0.750 4.710 0.920 ;
        RECT  4.250 0.275 4.340 1.295 ;
        RECT  3.960 0.425 4.250 0.595 ;
        RECT  3.900 1.185 4.250 1.295 ;
        RECT  3.865 0.905 3.975 1.015 ;
        RECT  3.775 0.275 3.865 1.015 ;
        RECT  3.565 0.275 3.775 0.365 ;
        RECT  3.595 0.465 3.685 1.505 ;
        RECT  3.515 0.465 3.595 0.575 ;
        RECT  3.555 1.085 3.595 1.505 ;
        RECT  3.395 0.255 3.565 0.365 ;
        RECT  3.335 0.455 3.425 1.295 ;
        RECT  2.825 0.275 3.395 0.365 ;
        RECT  3.290 0.455 3.335 0.645 ;
        RECT  3.295 1.085 3.335 1.295 ;
        RECT  3.020 1.085 3.295 1.185 ;
        RECT  3.200 0.735 3.245 0.905 ;
        RECT  3.110 0.485 3.200 0.905 ;
        RECT  2.785 0.485 3.110 0.575 ;
        RECT  2.915 0.710 3.020 1.185 ;
        RECT  2.655 0.255 2.825 0.365 ;
        RECT  2.695 0.485 2.785 1.185 ;
        RECT  2.540 0.485 2.695 0.595 ;
        RECT  2.665 1.075 2.695 1.185 ;
        RECT  2.555 1.075 2.665 1.430 ;
        RECT  2.370 0.780 2.495 0.890 ;
        RECT  2.060 1.395 2.440 1.510 ;
        RECT  2.250 0.255 2.420 0.405 ;
        RECT  2.275 0.525 2.370 1.135 ;
        RECT  2.040 0.525 2.275 0.635 ;
        RECT  2.065 1.025 2.275 1.135 ;
        RECT  0.865 0.305 2.250 0.405 ;
        RECT  1.950 0.800 2.115 0.910 ;
        RECT  1.970 1.295 2.060 1.510 ;
        RECT  0.945 1.295 1.970 1.385 ;
        RECT  1.860 0.495 1.950 1.195 ;
        RECT  1.545 0.495 1.860 0.605 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.260 0.500 1.360 0.845 ;
        RECT  0.850 0.500 1.260 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.500 0.850 0.915 ;
        RECT  0.355 0.500 0.740 0.590 ;
        RECT  0.265 0.500 0.355 1.290 ;
        RECT  0.185 0.500 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFND0

MACRO SDFND1
    CLASS CORE ;
    FOREIGN SDFND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.285 5.350 1.490 ;
        RECT  5.215 0.285 5.250 0.665 ;
        RECT  5.215 1.050 5.250 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.455 4.575 0.645 ;
        RECT  4.550 1.045 4.565 1.290 ;
        RECT  4.450 0.455 4.550 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.400 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.190 1.635 5.400 1.965 ;
        RECT  3.080 1.385 3.190 1.965 ;
        RECT  1.760 1.635 3.080 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.750 5.160 0.920 ;
        RECT  4.985 0.275 5.075 0.920 ;
        RECT  4.340 0.275 4.985 0.365 ;
        RECT  4.710 0.455 4.825 1.245 ;
        RECT  4.535 1.415 4.745 1.525 ;
        RECT  4.650 0.750 4.710 0.920 ;
        RECT  3.735 1.435 4.535 1.525 ;
        RECT  4.250 0.275 4.340 1.345 ;
        RECT  3.975 0.475 4.250 0.645 ;
        RECT  3.920 1.245 4.250 1.345 ;
        RECT  3.885 1.015 4.035 1.125 ;
        RECT  3.795 0.275 3.885 1.125 ;
        RECT  3.630 0.275 3.795 0.365 ;
        RECT  3.705 1.330 3.735 1.525 ;
        RECT  3.595 0.465 3.705 1.525 ;
        RECT  3.460 0.255 3.630 0.365 ;
        RECT  3.395 0.455 3.485 1.295 ;
        RECT  2.885 0.275 3.460 0.365 ;
        RECT  3.350 0.455 3.395 0.645 ;
        RECT  3.365 1.085 3.395 1.295 ;
        RECT  3.080 1.085 3.365 1.185 ;
        RECT  3.260 0.735 3.305 0.905 ;
        RECT  3.170 0.485 3.260 0.905 ;
        RECT  2.845 0.485 3.170 0.575 ;
        RECT  2.975 0.825 3.080 1.185 ;
        RECT  2.715 0.255 2.885 0.365 ;
        RECT  2.755 0.485 2.845 1.175 ;
        RECT  2.610 0.485 2.755 0.595 ;
        RECT  2.725 1.065 2.755 1.175 ;
        RECT  2.615 1.065 2.725 1.430 ;
        RECT  2.430 0.780 2.570 0.890 ;
        RECT  2.120 1.395 2.500 1.510 ;
        RECT  2.320 0.255 2.490 0.405 ;
        RECT  2.335 0.545 2.430 1.135 ;
        RECT  2.110 0.545 2.335 0.655 ;
        RECT  2.140 1.025 2.335 1.135 ;
        RECT  0.865 0.305 2.320 0.405 ;
        RECT  2.020 0.800 2.175 0.910 ;
        RECT  2.030 1.295 2.120 1.510 ;
        RECT  1.460 1.295 2.030 1.385 ;
        RECT  1.920 0.510 2.020 1.165 ;
        RECT  1.615 0.510 1.920 0.620 ;
        RECT  1.555 1.055 1.920 1.165 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFND1

MACRO SDFND2
    CLASS CORE ;
    FOREIGN SDFND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.565 5.750 1.150 ;
        RECT  5.645 0.565 5.650 0.665 ;
        RECT  5.645 1.050 5.650 1.150 ;
        RECT  5.535 0.285 5.645 0.665 ;
        RECT  5.535 1.050 5.645 1.460 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.350 1.180 4.665 1.290 ;
        RECT  4.350 0.510 4.615 0.690 ;
        RECT  4.250 0.510 4.350 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.905 -0.165 6.000 0.165 ;
        RECT  5.795 -0.165 5.905 0.475 ;
        RECT  0.520 -0.165 5.795 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.905 1.635 6.000 1.965 ;
        RECT  5.795 1.250 5.905 1.965 ;
        RECT  5.385 1.635 5.795 1.965 ;
        RECT  5.275 1.050 5.385 1.965 ;
        RECT  3.190 1.635 5.275 1.965 ;
        RECT  3.080 1.385 3.190 1.965 ;
        RECT  1.760 1.635 3.080 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.365 0.750 5.480 0.920 ;
        RECT  5.275 0.275 5.365 0.920 ;
        RECT  4.160 0.275 5.275 0.365 ;
        RECT  5.085 0.505 5.175 1.460 ;
        RECT  4.795 0.505 5.085 0.615 ;
        RECT  5.015 1.250 5.085 1.460 ;
        RECT  4.925 0.750 4.995 1.110 ;
        RECT  4.885 0.750 4.925 1.505 ;
        RECT  4.835 1.020 4.885 1.505 ;
        RECT  3.745 1.395 4.835 1.505 ;
        RECT  4.705 0.505 4.795 0.890 ;
        RECT  4.460 0.780 4.705 0.890 ;
        RECT  4.070 0.275 4.160 1.295 ;
        RECT  4.020 0.425 4.070 0.595 ;
        RECT  3.960 1.185 4.070 1.295 ;
        RECT  3.925 0.875 3.980 1.045 ;
        RECT  3.835 0.275 3.925 1.045 ;
        RECT  3.630 0.275 3.835 0.365 ;
        RECT  3.655 0.465 3.745 1.505 ;
        RECT  3.575 0.465 3.655 0.575 ;
        RECT  3.585 1.385 3.655 1.505 ;
        RECT  3.460 0.255 3.630 0.365 ;
        RECT  3.395 0.455 3.485 1.295 ;
        RECT  2.885 0.275 3.460 0.365 ;
        RECT  3.350 0.455 3.395 0.645 ;
        RECT  3.365 1.085 3.395 1.295 ;
        RECT  3.080 1.085 3.365 1.185 ;
        RECT  3.260 0.735 3.305 0.905 ;
        RECT  3.170 0.485 3.260 0.905 ;
        RECT  2.845 0.485 3.170 0.575 ;
        RECT  2.975 0.825 3.080 1.185 ;
        RECT  2.715 0.255 2.885 0.365 ;
        RECT  2.755 0.485 2.845 1.175 ;
        RECT  2.610 0.485 2.755 0.595 ;
        RECT  2.725 1.065 2.755 1.175 ;
        RECT  2.615 1.065 2.725 1.430 ;
        RECT  2.430 0.780 2.570 0.890 ;
        RECT  2.120 1.395 2.500 1.510 ;
        RECT  2.320 0.255 2.490 0.405 ;
        RECT  2.335 0.545 2.430 1.135 ;
        RECT  2.110 0.545 2.335 0.655 ;
        RECT  2.140 1.025 2.335 1.135 ;
        RECT  0.865 0.305 2.320 0.405 ;
        RECT  2.020 0.800 2.175 0.910 ;
        RECT  2.030 1.295 2.120 1.510 ;
        RECT  1.460 1.295 2.030 1.385 ;
        RECT  1.920 0.510 2.020 1.165 ;
        RECT  1.615 0.510 1.920 0.620 ;
        RECT  1.555 1.055 1.920 1.165 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFND2

MACRO SDFND4
    CLASS CORE ;
    FOREIGN SDFND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.325 7.150 0.635 ;
        RECT  7.050 1.100 7.150 1.405 ;
        RECT  6.750 0.325 7.050 1.405 ;
        RECT  6.435 0.325 6.750 0.635 ;
        RECT  6.435 1.100 6.750 1.405 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 1.100 6.150 1.410 ;
        RECT  6.050 0.520 6.105 0.690 ;
        RECT  5.750 0.520 6.050 1.410 ;
        RECT  5.435 0.520 5.750 0.690 ;
        RECT  5.435 1.100 5.750 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 7.400 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.635 7.400 1.965 ;
        RECT  3.070 1.385 3.180 1.965 ;
        RECT  0.470 1.635 3.070 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.435 0.325 6.650 0.635 ;
        RECT  6.435 1.100 6.650 1.405 ;
        RECT  5.435 0.520 5.650 0.690 ;
        RECT  5.435 1.100 5.650 1.410 ;
        RECT  6.315 0.780 6.500 0.890 ;
        RECT  6.215 0.315 6.315 0.890 ;
        RECT  4.200 0.315 6.215 0.405 ;
        RECT  5.135 0.780 5.500 0.890 ;
        RECT  5.045 0.515 5.135 1.410 ;
        RECT  4.580 0.515 5.045 0.625 ;
        RECT  4.915 1.300 5.045 1.410 ;
        RECT  4.845 0.750 4.955 1.190 ;
        RECT  4.805 1.080 4.845 1.190 ;
        RECT  4.695 1.080 4.805 1.525 ;
        RECT  3.715 1.420 4.695 1.525 ;
        RECT  4.200 1.220 4.605 1.330 ;
        RECT  4.470 0.515 4.580 0.930 ;
        RECT  4.100 0.315 4.200 1.330 ;
        RECT  3.985 0.475 4.100 0.645 ;
        RECT  3.895 1.220 4.100 1.330 ;
        RECT  3.895 0.755 3.995 1.095 ;
        RECT  3.885 0.275 3.895 1.095 ;
        RECT  3.805 0.275 3.885 0.845 ;
        RECT  3.625 0.275 3.805 0.365 ;
        RECT  3.615 0.455 3.715 1.525 ;
        RECT  3.455 0.255 3.625 0.365 ;
        RECT  3.605 0.455 3.615 0.665 ;
        RECT  3.395 0.455 3.485 1.295 ;
        RECT  2.885 0.275 3.455 0.365 ;
        RECT  3.350 0.455 3.395 0.645 ;
        RECT  3.355 1.085 3.395 1.295 ;
        RECT  3.080 1.085 3.355 1.185 ;
        RECT  3.260 0.735 3.305 0.905 ;
        RECT  3.170 0.485 3.260 0.905 ;
        RECT  2.845 0.485 3.170 0.575 ;
        RECT  2.975 0.710 3.080 1.185 ;
        RECT  2.715 0.255 2.885 0.365 ;
        RECT  2.755 0.485 2.845 1.175 ;
        RECT  2.600 0.485 2.755 0.595 ;
        RECT  2.725 1.065 2.755 1.175 ;
        RECT  2.615 1.065 2.725 1.430 ;
        RECT  2.430 0.780 2.560 0.890 ;
        RECT  2.315 1.385 2.500 1.525 ;
        RECT  2.310 0.255 2.480 0.405 ;
        RECT  2.335 0.545 2.430 1.175 ;
        RECT  2.110 0.545 2.335 0.655 ;
        RECT  2.090 1.065 2.335 1.175 ;
        RECT  0.945 1.435 2.315 1.525 ;
        RECT  0.865 0.305 2.310 0.405 ;
        RECT  2.000 0.800 2.175 0.910 ;
        RECT  1.900 0.510 2.000 1.325 ;
        RECT  1.615 0.510 1.900 0.620 ;
        RECT  1.565 1.215 1.900 1.325 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFND4

MACRO SDFNSND0
    CLASS CORE ;
    FOREIGN SDFNSND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.630 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.470 6.150 1.290 ;
        RECT  6.025 0.470 6.050 0.675 ;
        RECT  6.025 1.020 6.050 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.490 5.750 1.120 ;
        RECT  5.515 0.490 5.650 0.660 ;
        RECT  5.625 1.020 5.650 1.120 ;
        RECT  5.515 1.020 5.625 1.230 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0355 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  1.000 0.710 1.050 0.920 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 6.200 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.635 6.200 1.965 ;
        RECT  5.730 1.455 5.840 1.965 ;
        RECT  5.120 1.635 5.730 1.965 ;
        RECT  5.010 1.455 5.120 1.965 ;
        RECT  4.650 1.635 5.010 1.965 ;
        RECT  4.480 1.395 4.650 1.965 ;
        RECT  3.730 1.635 4.480 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  1.760 1.635 3.620 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.935 0.760 5.960 0.930 ;
        RECT  5.845 0.275 5.935 0.930 ;
        RECT  4.655 0.275 5.845 0.365 ;
        RECT  5.420 0.750 5.560 0.920 ;
        RECT  5.330 0.475 5.420 1.525 ;
        RECT  5.000 0.475 5.330 0.585 ;
        RECT  5.280 1.315 5.330 1.525 ;
        RECT  5.190 0.750 5.240 0.920 ;
        RECT  5.100 0.750 5.190 1.305 ;
        RECT  4.170 1.215 5.100 1.305 ;
        RECT  4.890 0.475 5.000 0.920 ;
        RECT  4.500 1.015 4.955 1.125 ;
        RECT  4.500 0.275 4.655 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  2.765 0.275 4.320 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  2.950 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.055 1.015 3.575 1.125 ;
        RECT  3.230 0.580 3.340 0.905 ;
        RECT  2.805 0.580 3.230 0.680 ;
        RECT  2.945 0.905 3.055 1.125 ;
        RECT  2.860 1.215 2.950 1.525 ;
        RECT  2.700 1.435 2.860 1.525 ;
        RECT  2.695 0.465 2.805 1.005 ;
        RECT  2.585 0.905 2.695 1.275 ;
        RECT  2.435 0.305 2.545 0.645 ;
        RECT  0.865 0.305 2.435 0.405 ;
        RECT  2.295 1.295 2.405 1.525 ;
        RECT  2.240 0.510 2.340 1.135 ;
        RECT  0.945 1.295 2.295 1.385 ;
        RECT  2.110 0.510 2.240 0.620 ;
        RECT  2.065 1.025 2.240 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.255 0.495 1.360 0.845 ;
        RECT  0.850 0.495 1.255 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.495 0.850 0.915 ;
        RECT  0.355 0.495 0.740 0.590 ;
        RECT  0.265 0.495 0.355 1.290 ;
        RECT  0.185 0.495 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNSND0

MACRO SDFNSND1
    CLASS CORE ;
    FOREIGN SDFNSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0823 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.275 6.150 1.490 ;
        RECT  6.025 0.275 6.050 0.675 ;
        RECT  6.015 1.050 6.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1380 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.490 5.750 1.120 ;
        RECT  5.515 0.490 5.650 0.660 ;
        RECT  5.625 1.020 5.650 1.120 ;
        RECT  5.515 1.020 5.625 1.260 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 6.200 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.660 1.635 6.200 1.965 ;
        RECT  4.490 1.395 4.660 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  1.760 1.635 3.620 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.935 0.760 5.960 0.930 ;
        RECT  5.845 0.275 5.935 0.930 ;
        RECT  4.655 0.275 5.845 0.365 ;
        RECT  5.420 0.750 5.560 0.920 ;
        RECT  5.330 0.475 5.420 1.525 ;
        RECT  5.000 0.475 5.330 0.585 ;
        RECT  5.305 1.315 5.330 1.525 ;
        RECT  5.190 0.750 5.240 0.920 ;
        RECT  5.100 0.750 5.190 1.305 ;
        RECT  4.170 1.215 5.100 1.305 ;
        RECT  4.890 0.475 5.000 0.920 ;
        RECT  4.500 1.015 4.965 1.125 ;
        RECT  4.500 0.275 4.655 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  2.765 0.275 4.320 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  2.950 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.055 1.015 3.575 1.125 ;
        RECT  3.230 0.580 3.340 0.905 ;
        RECT  2.805 0.580 3.230 0.680 ;
        RECT  2.945 0.905 3.055 1.125 ;
        RECT  2.860 1.215 2.950 1.525 ;
        RECT  2.700 1.435 2.860 1.525 ;
        RECT  2.695 0.465 2.805 1.005 ;
        RECT  2.585 0.905 2.695 1.275 ;
        RECT  2.435 0.305 2.545 0.645 ;
        RECT  0.865 0.305 2.435 0.405 ;
        RECT  2.295 1.295 2.405 1.525 ;
        RECT  2.240 0.510 2.340 1.135 ;
        RECT  1.460 1.295 2.295 1.385 ;
        RECT  2.110 0.510 2.240 0.620 ;
        RECT  2.065 1.025 2.240 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.165 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.055 1.860 1.165 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNSND1

MACRO SDFNSND2
    CLASS CORE ;
    FOREIGN SDFNSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.1093 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.625 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.575 6.550 1.150 ;
        RECT  6.445 0.575 6.450 0.675 ;
        RECT  6.445 1.050 6.450 1.150 ;
        RECT  6.335 0.275 6.445 0.675 ;
        RECT  6.335 1.050 6.445 1.460 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.490 5.950 1.490 ;
        RECT  5.815 0.490 5.850 0.660 ;
        RECT  5.815 1.020 5.850 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.705 -0.165 6.800 0.165 ;
        RECT  6.595 -0.165 6.705 0.480 ;
        RECT  0.520 -0.165 6.595 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.705 1.635 6.800 1.965 ;
        RECT  6.595 1.250 6.705 1.965 ;
        RECT  6.185 1.635 6.595 1.965 ;
        RECT  6.075 1.250 6.185 1.965 ;
        RECT  5.665 1.635 6.075 1.965 ;
        RECT  5.555 1.050 5.665 1.965 ;
        RECT  4.660 1.635 5.555 1.965 ;
        RECT  4.490 1.395 4.660 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  1.760 1.635 3.620 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.170 0.790 6.340 0.900 ;
        RECT  6.070 0.275 6.170 0.900 ;
        RECT  4.655 0.275 6.070 0.365 ;
        RECT  5.435 0.750 5.760 0.920 ;
        RECT  5.345 0.475 5.435 1.525 ;
        RECT  5.000 0.475 5.345 0.585 ;
        RECT  5.295 1.315 5.345 1.525 ;
        RECT  5.205 0.750 5.255 0.920 ;
        RECT  5.115 0.750 5.205 1.305 ;
        RECT  4.170 1.215 5.115 1.305 ;
        RECT  4.890 0.475 5.000 0.920 ;
        RECT  4.500 1.015 4.940 1.125 ;
        RECT  4.500 0.275 4.655 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  2.765 0.275 4.320 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  2.950 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.055 1.015 3.575 1.125 ;
        RECT  3.230 0.580 3.340 0.905 ;
        RECT  2.805 0.580 3.230 0.680 ;
        RECT  2.945 0.905 3.055 1.125 ;
        RECT  2.860 1.215 2.950 1.525 ;
        RECT  2.700 1.435 2.860 1.525 ;
        RECT  2.695 0.465 2.805 1.005 ;
        RECT  2.585 0.905 2.695 1.275 ;
        RECT  2.435 0.305 2.545 0.645 ;
        RECT  0.865 0.305 2.435 0.405 ;
        RECT  2.295 1.295 2.405 1.525 ;
        RECT  2.240 0.510 2.340 1.135 ;
        RECT  1.460 1.295 2.295 1.385 ;
        RECT  2.110 0.510 2.240 0.620 ;
        RECT  2.065 1.025 2.240 1.135 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.165 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.055 1.860 1.165 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNSND2

MACRO SDFNSND4
    CLASS CORE ;
    FOREIGN SDFNSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.1093 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.625 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.320 7.475 0.630 ;
        RECT  7.250 1.100 7.475 1.410 ;
        RECT  6.950 0.320 7.250 1.410 ;
        RECT  6.805 0.320 6.950 0.630 ;
        RECT  6.805 1.100 6.950 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.520 6.455 0.690 ;
        RECT  6.250 1.100 6.455 1.410 ;
        RECT  5.950 0.520 6.250 1.410 ;
        RECT  5.775 0.520 5.950 0.690 ;
        RECT  5.775 1.100 5.950 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 -0.165 7.800 0.165 ;
        RECT  7.595 -0.165 7.705 0.680 ;
        RECT  0.520 -0.165 7.595 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 1.635 7.800 1.965 ;
        RECT  7.595 1.050 7.705 1.965 ;
        RECT  6.685 1.635 7.595 1.965 ;
        RECT  6.575 1.050 6.685 1.965 ;
        RECT  5.655 1.635 6.575 1.965 ;
        RECT  5.545 1.050 5.655 1.965 ;
        RECT  4.660 1.635 5.545 1.965 ;
        RECT  4.490 1.395 4.660 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  0.470 1.635 3.620 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.380 0.320 7.475 0.630 ;
        RECT  7.380 1.100 7.475 1.410 ;
        RECT  6.805 0.320 6.850 0.630 ;
        RECT  6.805 1.100 6.850 1.410 ;
        RECT  6.350 0.520 6.455 0.690 ;
        RECT  6.350 1.100 6.455 1.410 ;
        RECT  5.775 0.520 5.850 0.690 ;
        RECT  5.775 1.100 5.850 1.410 ;
        RECT  6.665 0.790 6.840 0.900 ;
        RECT  6.575 0.275 6.665 0.900 ;
        RECT  4.655 0.275 6.575 0.365 ;
        RECT  5.425 0.780 5.790 0.890 ;
        RECT  5.335 0.475 5.425 1.525 ;
        RECT  5.000 0.475 5.335 0.585 ;
        RECT  5.285 1.315 5.335 1.525 ;
        RECT  5.195 0.750 5.245 0.920 ;
        RECT  5.105 0.750 5.195 1.305 ;
        RECT  4.170 1.215 5.105 1.305 ;
        RECT  4.890 0.475 5.000 0.920 ;
        RECT  4.520 1.015 4.940 1.125 ;
        RECT  4.520 0.275 4.655 0.405 ;
        RECT  4.430 0.275 4.520 1.125 ;
        RECT  4.085 0.545 4.430 0.655 ;
        RECT  4.275 1.015 4.430 1.125 ;
        RECT  2.775 0.275 4.340 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.965 0.835 4.070 0.925 ;
        RECT  3.855 0.495 3.965 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.705 1.015 3.940 1.125 ;
        RECT  2.950 1.215 3.855 1.305 ;
        RECT  3.595 0.495 3.705 1.125 ;
        RECT  3.060 1.015 3.595 1.125 ;
        RECT  3.240 0.580 3.350 0.905 ;
        RECT  2.805 0.580 3.240 0.680 ;
        RECT  2.945 0.905 3.060 1.125 ;
        RECT  2.860 1.215 2.950 1.525 ;
        RECT  2.700 1.435 2.860 1.525 ;
        RECT  2.695 0.465 2.805 1.005 ;
        RECT  2.585 0.905 2.695 1.275 ;
        RECT  2.435 0.305 2.545 0.645 ;
        RECT  0.865 0.305 2.435 0.405 ;
        RECT  2.295 1.295 2.405 1.525 ;
        RECT  2.225 0.510 2.335 1.145 ;
        RECT  0.945 1.435 2.295 1.525 ;
        RECT  2.110 0.510 2.225 0.620 ;
        RECT  2.065 1.035 2.225 1.145 ;
        RECT  1.960 0.780 2.115 0.890 ;
        RECT  1.860 0.510 1.960 1.325 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.215 1.860 1.325 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFNSND4

MACRO SDFQD0
    CLASS CORE ;
    FOREIGN SDFQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.710 0.570 1.110 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0602 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.170 1.110 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.650 0.275 4.750 1.500 ;
        RECT  4.615 0.275 4.650 0.445 ;
        RECT  4.615 1.290 4.650 1.500 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 0.925 ;
        RECT  0.965 0.740 1.050 0.925 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0221 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.670 1.550 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.340 -0.165 4.800 0.165 ;
        RECT  4.230 -0.165 4.340 0.345 ;
        RECT  2.180 -0.165 4.230 0.165 ;
        RECT  2.080 -0.165 2.180 0.685 ;
        RECT  0.470 -0.165 2.080 0.165 ;
        RECT  0.360 -0.165 0.470 0.415 ;
        RECT  0.000 -0.165 0.360 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.340 1.635 4.800 1.965 ;
        RECT  4.230 1.455 4.340 1.965 ;
        RECT  3.220 1.635 4.230 1.965 ;
        RECT  3.050 1.445 3.220 1.965 ;
        RECT  2.440 1.635 3.050 1.965 ;
        RECT  2.350 1.105 2.440 1.965 ;
        RECT  2.195 1.105 2.350 1.215 ;
        RECT  0.500 1.635 2.350 1.965 ;
        RECT  2.085 1.025 2.195 1.215 ;
        RECT  0.330 1.435 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.470 0.565 4.560 1.105 ;
        RECT  4.070 0.565 4.470 0.675 ;
        RECT  4.440 1.000 4.470 1.105 ;
        RECT  4.340 1.000 4.440 1.195 ;
        RECT  4.250 0.800 4.380 0.910 ;
        RECT  4.160 0.800 4.250 1.345 ;
        RECT  3.775 1.235 4.160 1.345 ;
        RECT  3.960 0.565 4.070 0.960 ;
        RECT  3.705 1.435 3.875 1.545 ;
        RECT  3.675 0.445 3.775 1.345 ;
        RECT  3.450 1.435 3.705 1.525 ;
        RECT  3.585 0.445 3.675 0.555 ;
        RECT  3.600 1.235 3.675 1.345 ;
        RECT  3.305 0.255 3.575 0.355 ;
        RECT  3.490 1.085 3.505 1.175 ;
        RECT  3.400 0.525 3.490 1.175 ;
        RECT  3.360 1.265 3.450 1.525 ;
        RECT  3.100 0.525 3.400 0.635 ;
        RECT  3.315 1.085 3.400 1.175 ;
        RECT  2.640 1.265 3.360 1.355 ;
        RECT  3.215 0.255 3.305 0.365 ;
        RECT  3.195 0.745 3.305 0.995 ;
        RECT  2.890 0.275 3.215 0.365 ;
        RECT  2.820 0.905 3.195 0.995 ;
        RECT  3.010 0.525 3.100 0.815 ;
        RECT  2.920 0.705 3.010 0.815 ;
        RECT  2.690 0.255 2.890 0.365 ;
        RECT  2.730 0.485 2.820 1.175 ;
        RECT  2.565 0.485 2.730 0.595 ;
        RECT  2.540 1.065 2.730 1.175 ;
        RECT  2.530 1.265 2.640 1.500 ;
        RECT  2.495 0.710 2.605 0.920 ;
        RECT  1.980 0.810 2.495 0.920 ;
        RECT  2.150 1.315 2.260 1.525 ;
        RECT  1.330 1.435 2.150 1.525 ;
        RECT  1.890 0.445 1.980 1.230 ;
        RECT  1.820 0.445 1.890 0.635 ;
        RECT  1.835 1.020 1.890 1.230 ;
        RECT  1.730 0.725 1.800 0.905 ;
        RECT  1.640 0.490 1.730 1.310 ;
        RECT  1.550 0.275 1.640 0.580 ;
        RECT  1.545 1.200 1.640 1.310 ;
        RECT  1.240 0.275 1.350 0.875 ;
        RECT  1.230 1.055 1.330 1.525 ;
        RECT  0.695 0.275 1.240 0.365 ;
        RECT  0.875 1.055 1.230 1.165 ;
        RECT  0.875 0.455 0.955 0.625 ;
        RECT  0.785 0.455 0.875 1.165 ;
        RECT  0.720 1.255 0.830 1.515 ;
        RECT  0.350 1.255 0.720 1.345 ;
        RECT  0.605 0.275 0.695 0.615 ;
        RECT  0.350 0.525 0.605 0.615 ;
        RECT  0.260 0.525 0.350 1.345 ;
        RECT  0.185 0.525 0.260 0.615 ;
        RECT  0.245 1.220 0.260 1.345 ;
        RECT  0.045 1.220 0.245 1.330 ;
        RECT  0.075 0.415 0.185 0.615 ;
    END
END SDFQD0

MACRO SDFQD1
    CLASS CORE ;
    FOREIGN SDFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.150 0.480 4.440 0.590 ;
        RECT  4.150 1.085 4.440 1.195 ;
        RECT  4.050 0.480 4.150 1.195 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.000 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.635 5.000 1.965 ;
        RECT  3.050 1.385 3.160 1.965 ;
        RECT  1.760 1.635 3.050 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.560 0.275 4.670 1.245 ;
        RECT  4.175 1.370 4.590 1.480 ;
        RECT  4.555 0.275 4.560 0.890 ;
        RECT  4.240 0.770 4.555 0.890 ;
        RECT  4.065 1.370 4.175 1.495 ;
        RECT  3.645 1.385 4.065 1.495 ;
        RECT  3.845 0.275 3.905 0.860 ;
        RECT  3.815 0.275 3.845 1.285 ;
        RECT  3.605 0.275 3.815 0.365 ;
        RECT  3.735 0.770 3.815 1.285 ;
        RECT  3.645 0.475 3.695 0.665 ;
        RECT  3.555 0.475 3.645 1.495 ;
        RECT  3.435 0.255 3.605 0.365 ;
        RECT  3.375 0.455 3.465 1.295 ;
        RECT  2.895 0.275 3.435 0.365 ;
        RECT  3.330 0.455 3.375 0.645 ;
        RECT  3.335 1.085 3.375 1.295 ;
        RECT  3.060 1.085 3.335 1.185 ;
        RECT  3.240 0.735 3.285 0.905 ;
        RECT  3.150 0.475 3.240 0.905 ;
        RECT  2.795 0.475 3.150 0.565 ;
        RECT  2.955 0.710 3.060 1.185 ;
        RECT  2.685 0.255 2.895 0.365 ;
        RECT  2.695 0.475 2.795 1.185 ;
        RECT  2.585 0.475 2.695 0.575 ;
        RECT  2.590 1.075 2.695 1.185 ;
        RECT  2.410 0.745 2.555 0.865 ;
        RECT  2.300 1.235 2.505 1.385 ;
        RECT  2.275 0.255 2.445 0.405 ;
        RECT  2.315 0.565 2.410 1.135 ;
        RECT  2.110 0.565 2.315 0.675 ;
        RECT  2.065 1.025 2.315 1.135 ;
        RECT  1.460 1.295 2.300 1.385 ;
        RECT  0.865 0.305 2.275 0.405 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFQD1

MACRO SDFQD2
    CLASS CORE ;
    FOREIGN SDFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.265 0.275 4.375 0.675 ;
        RECT  4.150 1.110 4.375 1.290 ;
        RECT  4.150 0.575 4.265 0.675 ;
        RECT  4.050 0.575 4.150 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.200 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.635 5.200 1.965 ;
        RECT  3.010 1.385 3.120 1.965 ;
        RECT  1.760 1.635 3.010 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.875 0.555 4.935 1.410 ;
        RECT  4.845 0.275 4.875 1.410 ;
        RECT  4.765 0.275 4.845 0.655 ;
        RECT  4.715 1.300 4.845 1.410 ;
        RECT  4.555 0.555 4.765 0.655 ;
        RECT  4.645 0.750 4.755 1.140 ;
        RECT  4.615 1.050 4.645 1.140 ;
        RECT  4.525 1.050 4.615 1.495 ;
        RECT  4.465 0.555 4.555 0.890 ;
        RECT  3.605 1.385 4.525 1.495 ;
        RECT  4.260 0.770 4.465 0.890 ;
        RECT  3.800 0.275 3.865 1.055 ;
        RECT  3.775 0.275 3.800 1.265 ;
        RECT  3.565 0.275 3.775 0.365 ;
        RECT  3.695 0.965 3.775 1.265 ;
        RECT  3.605 0.465 3.655 0.665 ;
        RECT  3.515 0.465 3.605 1.495 ;
        RECT  3.395 0.255 3.565 0.365 ;
        RECT  3.335 0.455 3.425 1.295 ;
        RECT  2.835 0.275 3.395 0.365 ;
        RECT  3.290 0.455 3.335 0.645 ;
        RECT  3.295 1.085 3.335 1.295 ;
        RECT  3.020 1.085 3.295 1.185 ;
        RECT  3.200 0.735 3.245 0.905 ;
        RECT  3.110 0.475 3.200 0.905 ;
        RECT  2.785 0.475 3.110 0.565 ;
        RECT  2.915 0.710 3.020 1.185 ;
        RECT  2.665 0.255 2.835 0.365 ;
        RECT  2.695 0.475 2.785 1.185 ;
        RECT  2.545 0.475 2.695 0.575 ;
        RECT  2.550 1.075 2.695 1.185 ;
        RECT  2.370 0.725 2.515 0.835 ;
        RECT  2.260 1.235 2.465 1.385 ;
        RECT  2.235 0.255 2.405 0.405 ;
        RECT  2.275 0.565 2.370 1.135 ;
        RECT  2.110 0.565 2.275 0.675 ;
        RECT  2.055 1.025 2.275 1.135 ;
        RECT  1.460 1.295 2.260 1.385 ;
        RECT  0.865 0.305 2.235 0.405 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFQD2

MACRO SDFQD4
    CLASS CORE ;
    FOREIGN SDFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.315 5.005 0.635 ;
        RECT  4.850 1.120 5.005 1.290 ;
        RECT  4.550 0.315 4.850 1.290 ;
        RECT  4.320 0.315 4.550 0.635 ;
        RECT  4.335 1.120 4.550 1.290 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 5.800 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.220 1.635 5.800 1.965 ;
        RECT  3.110 1.385 3.220 1.965 ;
        RECT  0.470 1.635 3.110 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.950 0.315 5.005 0.635 ;
        RECT  4.950 1.120 5.005 1.290 ;
        RECT  4.320 0.315 4.450 0.635 ;
        RECT  4.335 1.120 4.450 1.290 ;
        RECT  5.560 0.555 5.650 1.410 ;
        RECT  5.475 0.555 5.560 0.655 ;
        RECT  5.315 1.300 5.560 1.410 ;
        RECT  5.365 0.275 5.475 0.655 ;
        RECT  5.360 0.750 5.470 1.140 ;
        RECT  5.215 0.555 5.365 0.655 ;
        RECT  5.215 1.050 5.360 1.140 ;
        RECT  5.125 0.555 5.215 0.890 ;
        RECT  5.125 1.050 5.215 1.495 ;
        RECT  4.970 0.780 5.125 0.890 ;
        RECT  3.705 1.385 5.125 1.495 ;
        RECT  3.900 0.275 3.965 1.055 ;
        RECT  3.875 0.275 3.900 1.265 ;
        RECT  3.665 0.275 3.875 0.365 ;
        RECT  3.795 0.965 3.875 1.265 ;
        RECT  3.705 0.465 3.755 0.665 ;
        RECT  3.615 0.465 3.705 1.495 ;
        RECT  3.495 0.255 3.665 0.365 ;
        RECT  3.435 0.455 3.525 1.295 ;
        RECT  2.935 0.275 3.495 0.365 ;
        RECT  3.390 0.455 3.435 0.645 ;
        RECT  3.395 1.085 3.435 1.295 ;
        RECT  3.120 1.085 3.395 1.185 ;
        RECT  3.300 0.735 3.345 0.905 ;
        RECT  3.210 0.475 3.300 0.905 ;
        RECT  2.885 0.475 3.210 0.565 ;
        RECT  3.015 0.710 3.120 1.185 ;
        RECT  2.765 0.255 2.935 0.365 ;
        RECT  2.795 0.475 2.885 1.185 ;
        RECT  2.645 0.475 2.795 0.575 ;
        RECT  2.650 1.075 2.795 1.185 ;
        RECT  2.470 0.745 2.615 0.855 ;
        RECT  2.360 1.240 2.565 1.385 ;
        RECT  0.865 0.305 2.520 0.405 ;
        RECT  2.375 0.545 2.470 1.135 ;
        RECT  2.110 0.545 2.375 0.655 ;
        RECT  2.080 1.025 2.375 1.135 ;
        RECT  1.460 1.295 2.360 1.385 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFQD4

MACRO SDFQND0
    CLASS CORE ;
    FOREIGN SDFQND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0498 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNAGATEAREA 0.0180 ;
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.260 0.275 4.350 1.490 ;
        RECT  4.200 0.275 4.260 0.640 ;
        RECT  4.050 1.310 4.260 1.490 ;
        RECT  3.950 0.530 4.200 0.640 ;
        RECT  3.850 0.530 3.950 0.920 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0354 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.100 ;
        RECT  1.000 0.710 1.050 0.880 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 4.400 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 1.635 4.400 1.965 ;
        RECT  2.960 1.385 3.070 1.965 ;
        RECT  1.730 1.635 2.960 1.965 ;
        RECT  1.540 1.495 1.730 1.965 ;
        RECT  0.470 1.635 1.540 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.060 0.730 4.170 1.145 ;
        RECT  3.950 1.045 4.060 1.145 ;
        RECT  3.860 1.045 3.950 1.495 ;
        RECT  3.550 1.385 3.860 1.495 ;
        RECT  3.670 0.275 3.760 1.285 ;
        RECT  3.515 0.275 3.670 0.365 ;
        RECT  3.645 1.095 3.670 1.285 ;
        RECT  3.550 0.475 3.580 0.645 ;
        RECT  3.460 0.475 3.550 1.495 ;
        RECT  3.345 0.255 3.515 0.365 ;
        RECT  3.280 0.455 3.370 1.295 ;
        RECT  2.785 0.275 3.345 0.365 ;
        RECT  3.230 0.455 3.280 0.645 ;
        RECT  3.245 1.085 3.280 1.295 ;
        RECT  2.960 1.085 3.245 1.185 ;
        RECT  3.140 0.735 3.190 0.905 ;
        RECT  3.050 0.475 3.140 0.905 ;
        RECT  2.735 0.475 3.050 0.565 ;
        RECT  2.860 0.710 2.960 1.185 ;
        RECT  2.615 0.255 2.785 0.365 ;
        RECT  2.645 0.475 2.735 1.185 ;
        RECT  2.495 0.475 2.645 0.575 ;
        RECT  2.495 1.075 2.645 1.185 ;
        RECT  2.335 0.735 2.460 0.845 ;
        RECT  2.235 1.235 2.410 1.385 ;
        RECT  2.185 0.255 2.355 0.405 ;
        RECT  2.240 0.565 2.335 1.115 ;
        RECT  2.045 0.565 2.240 0.675 ;
        RECT  2.140 1.005 2.240 1.115 ;
        RECT  0.945 1.295 2.235 1.385 ;
        RECT  0.865 0.305 2.185 0.405 ;
        RECT  2.025 1.005 2.140 1.195 ;
        RECT  1.930 0.800 2.080 0.910 ;
        RECT  1.840 0.495 1.930 1.195 ;
        RECT  1.550 0.495 1.840 0.605 ;
        RECT  1.525 1.085 1.840 1.195 ;
        RECT  1.240 0.500 1.350 0.865 ;
        RECT  0.850 0.500 1.240 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.500 0.850 0.915 ;
        RECT  0.355 0.500 0.740 0.590 ;
        RECT  0.265 0.500 0.355 1.290 ;
        RECT  0.185 0.500 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFQND0

MACRO SDFQND1
    CLASS CORE ;
    FOREIGN SDFQND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.815 0.275 4.950 1.490 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.640 -0.165 5.000 0.165 ;
        RECT  4.530 -0.165 4.640 0.345 ;
        RECT  4.155 -0.165 4.530 0.165 ;
        RECT  4.045 -0.165 4.155 0.345 ;
        RECT  0.520 -0.165 4.045 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.635 5.000 1.965 ;
        RECT  3.020 1.385 3.130 1.965 ;
        RECT  1.760 1.635 3.020 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.605 0.505 4.705 1.495 ;
        RECT  4.035 0.505 4.605 0.615 ;
        RECT  4.295 1.385 4.605 1.495 ;
        RECT  4.385 0.730 4.495 1.255 ;
        RECT  4.140 1.150 4.385 1.255 ;
        RECT  4.040 1.150 4.140 1.495 ;
        RECT  3.635 1.385 4.040 1.495 ;
        RECT  3.925 0.505 4.035 0.940 ;
        RECT  3.745 0.275 3.835 1.290 ;
        RECT  3.575 0.275 3.745 0.365 ;
        RECT  3.725 1.120 3.745 1.290 ;
        RECT  3.635 0.455 3.655 0.665 ;
        RECT  3.545 0.455 3.635 1.495 ;
        RECT  3.405 0.255 3.575 0.365 ;
        RECT  3.515 1.385 3.545 1.495 ;
        RECT  3.345 0.455 3.435 1.295 ;
        RECT  2.845 0.275 3.405 0.365 ;
        RECT  3.300 0.455 3.345 0.645 ;
        RECT  3.305 1.085 3.345 1.295 ;
        RECT  3.030 1.085 3.305 1.185 ;
        RECT  3.210 0.735 3.255 0.905 ;
        RECT  3.120 0.475 3.210 0.905 ;
        RECT  2.795 0.475 3.120 0.565 ;
        RECT  2.925 0.710 3.030 1.185 ;
        RECT  2.675 0.255 2.845 0.365 ;
        RECT  2.705 0.475 2.795 1.185 ;
        RECT  2.555 0.475 2.705 0.575 ;
        RECT  2.560 1.075 2.705 1.185 ;
        RECT  2.380 0.735 2.525 0.845 ;
        RECT  2.270 1.235 2.475 1.385 ;
        RECT  2.245 0.255 2.415 0.405 ;
        RECT  2.275 0.565 2.380 1.135 ;
        RECT  2.110 0.565 2.275 0.675 ;
        RECT  2.065 1.025 2.275 1.135 ;
        RECT  1.460 1.295 2.270 1.385 ;
        RECT  0.865 0.305 2.245 0.405 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFQND1

MACRO SDFQND2
    CLASS CORE ;
    FOREIGN SDFQND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.285 4.950 1.490 ;
        RECT  4.765 0.285 4.850 0.665 ;
        RECT  4.765 1.050 4.850 1.490 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.590 -0.165 5.200 0.165 ;
        RECT  4.480 -0.165 4.590 0.345 ;
        RECT  0.520 -0.165 4.480 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.125 1.635 5.200 1.965 ;
        RECT  3.015 1.385 3.125 1.965 ;
        RECT  1.760 1.635 3.015 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.585 0.505 4.675 1.495 ;
        RECT  4.045 0.505 4.585 0.615 ;
        RECT  4.220 1.385 4.585 1.495 ;
        RECT  4.345 0.740 4.455 1.235 ;
        RECT  4.110 1.145 4.345 1.235 ;
        RECT  4.020 1.145 4.110 1.495 ;
        RECT  3.935 0.505 4.045 0.940 ;
        RECT  3.610 1.385 4.020 1.495 ;
        RECT  3.800 0.275 3.840 0.845 ;
        RECT  3.750 0.275 3.800 1.275 ;
        RECT  3.570 0.275 3.750 0.365 ;
        RECT  3.700 0.755 3.750 1.275 ;
        RECT  3.610 0.465 3.660 0.645 ;
        RECT  3.520 0.465 3.610 1.495 ;
        RECT  3.400 0.255 3.570 0.365 ;
        RECT  3.340 0.455 3.430 1.295 ;
        RECT  2.845 0.275 3.400 0.365 ;
        RECT  3.295 0.455 3.340 0.645 ;
        RECT  3.300 1.085 3.340 1.295 ;
        RECT  3.025 1.085 3.300 1.185 ;
        RECT  3.205 0.735 3.250 0.905 ;
        RECT  3.115 0.475 3.205 0.905 ;
        RECT  2.795 0.475 3.115 0.565 ;
        RECT  2.920 0.685 3.025 1.185 ;
        RECT  2.675 0.255 2.845 0.365 ;
        RECT  2.705 0.475 2.795 1.185 ;
        RECT  2.555 0.475 2.705 0.575 ;
        RECT  2.555 1.075 2.705 1.185 ;
        RECT  2.380 0.735 2.525 0.845 ;
        RECT  2.265 1.235 2.470 1.385 ;
        RECT  2.245 0.255 2.415 0.405 ;
        RECT  2.285 0.565 2.380 1.135 ;
        RECT  2.110 0.565 2.285 0.675 ;
        RECT  2.060 1.025 2.285 1.135 ;
        RECT  1.460 1.295 2.265 1.385 ;
        RECT  0.865 0.305 2.245 0.405 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFQND2

MACRO SDFQND4
    CLASS CORE ;
    FOREIGN SDFQND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.325 5.475 0.635 ;
        RECT  5.250 1.155 5.475 1.465 ;
        RECT  4.950 0.325 5.250 1.465 ;
        RECT  4.805 0.325 4.950 0.635 ;
        RECT  4.805 1.155 4.950 1.465 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.705 -0.165 5.800 0.165 ;
        RECT  5.595 -0.165 5.705 0.685 ;
        RECT  4.660 -0.165 5.595 0.165 ;
        RECT  4.550 -0.165 4.660 0.345 ;
        RECT  0.520 -0.165 4.550 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.705 1.635 5.800 1.965 ;
        RECT  5.595 1.105 5.705 1.965 ;
        RECT  3.195 1.635 5.595 1.965 ;
        RECT  3.085 1.385 3.195 1.965 ;
        RECT  0.470 1.635 3.085 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.350 0.325 5.475 0.635 ;
        RECT  5.350 1.155 5.475 1.465 ;
        RECT  4.805 0.325 4.850 0.635 ;
        RECT  4.805 1.155 4.850 1.465 ;
        RECT  4.595 0.505 4.695 1.495 ;
        RECT  4.115 0.505 4.595 0.615 ;
        RECT  4.290 1.385 4.595 1.495 ;
        RECT  4.375 0.740 4.485 1.235 ;
        RECT  4.180 1.145 4.375 1.235 ;
        RECT  4.090 1.145 4.180 1.495 ;
        RECT  4.005 0.505 4.115 0.940 ;
        RECT  3.680 1.385 4.090 1.495 ;
        RECT  3.870 0.275 3.910 0.845 ;
        RECT  3.820 0.275 3.870 1.275 ;
        RECT  3.640 0.275 3.820 0.365 ;
        RECT  3.770 0.755 3.820 1.275 ;
        RECT  3.680 0.465 3.730 0.645 ;
        RECT  3.590 0.465 3.680 1.495 ;
        RECT  3.470 0.255 3.640 0.365 ;
        RECT  3.410 0.455 3.500 1.295 ;
        RECT  2.915 0.275 3.470 0.365 ;
        RECT  3.365 0.455 3.410 0.645 ;
        RECT  3.370 1.085 3.410 1.295 ;
        RECT  3.095 1.085 3.370 1.185 ;
        RECT  3.275 0.735 3.320 0.905 ;
        RECT  3.185 0.475 3.275 0.905 ;
        RECT  2.865 0.475 3.185 0.565 ;
        RECT  2.990 0.685 3.095 1.185 ;
        RECT  2.745 0.255 2.915 0.365 ;
        RECT  2.775 0.475 2.865 1.185 ;
        RECT  2.625 0.475 2.775 0.575 ;
        RECT  2.625 1.075 2.775 1.185 ;
        RECT  2.450 0.735 2.595 0.845 ;
        RECT  2.335 1.235 2.540 1.385 ;
        RECT  0.865 0.305 2.510 0.405 ;
        RECT  2.355 0.545 2.450 1.135 ;
        RECT  2.110 0.545 2.355 0.655 ;
        RECT  2.080 1.025 2.355 1.135 ;
        RECT  1.460 1.295 2.335 1.385 ;
        RECT  1.960 0.800 2.115 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFQND4

MACRO SDFSND0
    CLASS CORE ;
    FOREIGN SDFSND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.470 6.150 1.290 ;
        RECT  6.025 0.470 6.050 0.675 ;
        RECT  6.025 1.020 6.050 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.490 5.750 1.120 ;
        RECT  5.515 0.490 5.650 0.660 ;
        RECT  5.625 1.020 5.650 1.120 ;
        RECT  5.515 1.020 5.625 1.230 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0355 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  1.000 0.710 1.050 0.920 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 6.200 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.635 6.200 1.965 ;
        RECT  5.730 1.455 5.840 1.965 ;
        RECT  5.130 1.635 5.730 1.965 ;
        RECT  5.020 1.455 5.130 1.965 ;
        RECT  4.660 1.635 5.020 1.965 ;
        RECT  4.490 1.395 4.660 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  1.760 1.635 3.620 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.935 0.760 5.960 0.930 ;
        RECT  5.845 0.275 5.935 0.930 ;
        RECT  4.655 0.275 5.845 0.365 ;
        RECT  5.420 0.750 5.560 0.920 ;
        RECT  5.330 0.475 5.420 1.525 ;
        RECT  5.000 0.475 5.330 0.585 ;
        RECT  5.280 1.315 5.330 1.525 ;
        RECT  5.190 0.750 5.240 0.920 ;
        RECT  5.100 0.750 5.190 1.305 ;
        RECT  4.170 1.215 5.100 1.305 ;
        RECT  4.890 0.475 5.000 0.920 ;
        RECT  4.500 1.015 4.965 1.125 ;
        RECT  4.500 0.275 4.655 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  3.105 0.275 4.320 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  3.335 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.045 1.015 3.575 1.125 ;
        RECT  3.230 0.495 3.340 0.905 ;
        RECT  3.245 1.215 3.335 1.525 ;
        RECT  2.635 1.425 3.245 1.525 ;
        RECT  2.700 0.495 3.230 0.605 ;
        RECT  2.745 0.275 3.105 0.365 ;
        RECT  2.935 0.900 3.045 1.125 ;
        RECT  2.590 0.495 2.700 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.275 1.295 2.445 1.445 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.080 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  0.945 1.295 2.275 1.385 ;
        RECT  1.960 0.780 2.135 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.255 0.495 1.360 0.845 ;
        RECT  0.850 0.495 1.255 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.495 0.850 0.915 ;
        RECT  0.355 0.495 0.740 0.590 ;
        RECT  0.265 0.495 0.355 1.290 ;
        RECT  0.185 0.495 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSND0

MACRO SDFSND1
    CLASS CORE ;
    FOREIGN SDFSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0823 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.275 6.150 1.490 ;
        RECT  6.025 0.275 6.050 0.675 ;
        RECT  6.015 1.050 6.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1380 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.490 5.750 1.120 ;
        RECT  5.515 0.490 5.650 0.660 ;
        RECT  5.625 1.020 5.650 1.120 ;
        RECT  5.515 1.020 5.625 1.260 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 6.200 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.660 1.635 6.200 1.965 ;
        RECT  4.490 1.395 4.660 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  3.215 1.635 3.620 1.965 ;
        RECT  3.045 1.395 3.215 1.965 ;
        RECT  1.760 1.635 3.045 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.935 0.760 5.960 0.930 ;
        RECT  5.845 0.275 5.935 0.930 ;
        RECT  4.655 0.275 5.845 0.365 ;
        RECT  5.420 0.750 5.560 0.920 ;
        RECT  5.330 0.475 5.420 1.525 ;
        RECT  5.000 0.475 5.330 0.585 ;
        RECT  5.305 1.315 5.330 1.525 ;
        RECT  5.190 0.750 5.240 0.920 ;
        RECT  5.100 0.750 5.190 1.305 ;
        RECT  4.170 1.215 5.100 1.305 ;
        RECT  4.890 0.475 5.000 0.920 ;
        RECT  4.500 1.015 4.965 1.125 ;
        RECT  4.500 0.275 4.655 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  2.745 0.275 4.320 0.385 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  2.930 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.045 1.015 3.575 1.125 ;
        RECT  3.230 0.495 3.340 0.905 ;
        RECT  2.700 0.495 3.230 0.605 ;
        RECT  2.935 0.900 3.045 1.125 ;
        RECT  2.840 1.215 2.930 1.525 ;
        RECT  2.635 1.425 2.840 1.525 ;
        RECT  2.590 0.495 2.700 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.275 1.295 2.445 1.445 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.080 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  1.460 1.295 2.275 1.385 ;
        RECT  1.960 0.780 2.135 0.890 ;
        RECT  1.860 0.510 1.960 1.165 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.055 1.860 1.165 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSND1

MACRO SDFSND2
    CLASS CORE ;
    FOREIGN SDFSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0823 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.630 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.575 6.550 1.150 ;
        RECT  6.445 0.575 6.450 0.675 ;
        RECT  6.445 1.050 6.450 1.150 ;
        RECT  6.335 0.285 6.445 0.675 ;
        RECT  6.335 1.050 6.445 1.460 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.475 5.950 1.490 ;
        RECT  5.815 0.475 5.850 0.675 ;
        RECT  5.815 1.020 5.850 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.705 -0.165 6.800 0.165 ;
        RECT  6.595 -0.165 6.705 0.475 ;
        RECT  0.520 -0.165 6.595 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.705 1.635 6.800 1.965 ;
        RECT  6.595 1.250 6.705 1.965 ;
        RECT  6.185 1.635 6.595 1.965 ;
        RECT  6.075 1.050 6.185 1.965 ;
        RECT  5.140 1.635 6.075 1.965 ;
        RECT  5.030 1.455 5.140 1.965 ;
        RECT  4.695 1.635 5.030 1.965 ;
        RECT  4.490 1.395 4.695 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  3.215 1.635 3.620 1.965 ;
        RECT  3.045 1.395 3.215 1.965 ;
        RECT  1.760 1.635 3.045 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.245 0.790 6.360 0.900 ;
        RECT  6.155 0.275 6.245 0.900 ;
        RECT  4.685 0.275 6.155 0.365 ;
        RECT  5.705 0.760 5.750 0.930 ;
        RECT  5.615 0.475 5.705 1.160 ;
        RECT  5.035 0.475 5.615 0.585 ;
        RECT  5.425 1.050 5.615 1.160 ;
        RECT  5.225 0.780 5.440 0.890 ;
        RECT  5.315 1.050 5.425 1.460 ;
        RECT  5.135 0.780 5.225 1.305 ;
        RECT  4.170 1.215 5.135 1.305 ;
        RECT  4.925 0.475 5.035 0.920 ;
        RECT  4.500 1.015 4.975 1.125 ;
        RECT  4.500 0.275 4.685 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  2.745 0.275 4.320 0.385 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  2.930 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.045 1.015 3.575 1.125 ;
        RECT  3.230 0.495 3.340 0.905 ;
        RECT  2.700 0.495 3.230 0.605 ;
        RECT  2.935 0.900 3.045 1.125 ;
        RECT  2.840 1.215 2.930 1.525 ;
        RECT  2.635 1.425 2.840 1.525 ;
        RECT  2.590 0.495 2.700 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.275 1.295 2.445 1.445 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.080 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  1.460 1.295 2.275 1.385 ;
        RECT  1.960 0.780 2.135 0.890 ;
        RECT  1.860 0.510 1.960 1.165 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.055 1.860 1.165 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSND2

MACRO SDFSND4
    CLASS CORE ;
    FOREIGN SDFSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.1093 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.630 0.510 4.750 0.925 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.325 7.475 0.635 ;
        RECT  7.250 1.100 7.475 1.410 ;
        RECT  6.950 0.325 7.250 1.410 ;
        RECT  6.795 0.325 6.950 0.635 ;
        RECT  6.795 1.100 6.950 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.525 6.445 0.690 ;
        RECT  6.250 1.100 6.445 1.410 ;
        RECT  5.950 0.525 6.250 1.410 ;
        RECT  5.775 0.525 5.950 0.695 ;
        RECT  5.775 1.100 5.950 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 -0.165 7.800 0.165 ;
        RECT  7.595 -0.165 7.705 0.685 ;
        RECT  0.520 -0.165 7.595 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 1.635 7.800 1.965 ;
        RECT  7.595 1.050 7.705 1.965 ;
        RECT  6.675 1.635 7.595 1.965 ;
        RECT  6.565 1.050 6.675 1.965 ;
        RECT  5.655 1.635 6.565 1.965 ;
        RECT  5.545 1.050 5.655 1.965 ;
        RECT  4.690 1.635 5.545 1.965 ;
        RECT  4.490 1.395 4.690 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  3.215 1.635 3.620 1.965 ;
        RECT  3.045 1.395 3.215 1.965 ;
        RECT  0.470 1.635 3.045 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.350 0.325 7.475 0.635 ;
        RECT  7.350 1.100 7.475 1.410 ;
        RECT  6.795 0.325 6.850 0.635 ;
        RECT  6.795 1.100 6.850 1.410 ;
        RECT  6.350 0.525 6.445 0.690 ;
        RECT  6.350 1.100 6.445 1.410 ;
        RECT  5.775 0.525 5.850 0.695 ;
        RECT  5.775 1.100 5.850 1.410 ;
        RECT  6.665 0.790 6.830 0.900 ;
        RECT  6.575 0.275 6.665 0.900 ;
        RECT  4.685 0.275 6.575 0.365 ;
        RECT  5.435 0.785 5.830 0.890 ;
        RECT  5.345 0.475 5.435 1.460 ;
        RECT  5.015 0.475 5.345 0.585 ;
        RECT  5.285 1.050 5.345 1.460 ;
        RECT  5.195 0.750 5.255 0.920 ;
        RECT  5.105 0.750 5.195 1.305 ;
        RECT  4.170 1.215 5.105 1.305 ;
        RECT  4.905 0.475 5.015 0.920 ;
        RECT  4.500 1.015 4.945 1.125 ;
        RECT  4.500 0.275 4.685 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  2.745 0.275 4.320 0.385 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  2.930 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.045 1.015 3.575 1.125 ;
        RECT  3.230 0.495 3.340 0.905 ;
        RECT  2.700 0.495 3.230 0.605 ;
        RECT  2.935 0.900 3.045 1.125 ;
        RECT  2.840 1.215 2.930 1.525 ;
        RECT  2.635 1.425 2.840 1.525 ;
        RECT  2.590 0.495 2.700 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.275 1.295 2.445 1.445 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.080 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  1.460 1.295 2.275 1.385 ;
        RECT  1.960 0.780 2.135 0.890 ;
        RECT  1.860 0.510 1.960 1.165 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.055 1.860 1.165 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSND4

MACRO SDFSNQD0
    CLASS CORE ;
    FOREIGN SDFSNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0790 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.510 4.750 0.925 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.520 5.950 1.180 ;
        RECT  5.525 0.520 5.850 0.630 ;
        RECT  5.525 1.070 5.850 1.180 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0355 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.710 1.150 1.090 ;
        RECT  1.000 0.710 1.050 0.920 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0217 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.165 6.000 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.890 1.635 6.000 1.965 ;
        RECT  5.780 1.455 5.890 1.965 ;
        RECT  5.130 1.635 5.780 1.965 ;
        RECT  5.020 1.455 5.130 1.965 ;
        RECT  4.660 1.635 5.020 1.965 ;
        RECT  4.490 1.395 4.660 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  1.760 1.635 3.620 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.430 0.780 5.760 0.890 ;
        RECT  5.340 0.330 5.430 1.265 ;
        RECT  5.000 0.330 5.340 0.440 ;
        RECT  5.305 1.055 5.340 1.265 ;
        RECT  5.190 0.750 5.250 0.920 ;
        RECT  5.100 0.750 5.190 1.305 ;
        RECT  4.170 1.215 5.100 1.305 ;
        RECT  4.890 0.330 5.000 0.920 ;
        RECT  4.500 1.015 4.965 1.125 ;
        RECT  4.500 0.275 4.655 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  3.105 0.275 4.320 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  3.335 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.045 1.015 3.575 1.125 ;
        RECT  3.230 0.495 3.340 0.905 ;
        RECT  3.245 1.215 3.335 1.525 ;
        RECT  2.635 1.425 3.245 1.525 ;
        RECT  2.700 0.495 3.230 0.605 ;
        RECT  2.745 0.275 3.105 0.365 ;
        RECT  2.935 0.900 3.045 1.125 ;
        RECT  2.590 0.495 2.700 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.275 1.295 2.445 1.445 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.080 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  0.945 1.295 2.275 1.385 ;
        RECT  1.960 0.780 2.135 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.255 0.495 1.360 0.845 ;
        RECT  0.850 0.495 1.255 0.590 ;
        RECT  0.835 1.145 0.945 1.385 ;
        RECT  0.740 0.495 0.850 0.915 ;
        RECT  0.355 0.495 0.740 0.590 ;
        RECT  0.265 0.495 0.355 1.290 ;
        RECT  0.185 0.495 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSNQD0

MACRO SDFSNQD1
    CLASS CORE ;
    FOREIGN SDFSNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0790 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.625 0.510 4.750 0.925 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.285 5.950 1.490 ;
        RECT  5.815 0.285 5.850 0.675 ;
        RECT  5.815 1.050 5.850 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.665 -0.165 6.000 0.165 ;
        RECT  5.555 -0.165 5.665 0.665 ;
        RECT  5.095 -0.165 5.555 0.165 ;
        RECT  4.985 -0.165 5.095 0.465 ;
        RECT  0.520 -0.165 4.985 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.665 1.635 6.000 1.965 ;
        RECT  5.555 1.070 5.665 1.965 ;
        RECT  4.660 1.635 5.555 1.965 ;
        RECT  4.490 1.395 4.660 1.965 ;
        RECT  3.730 1.635 4.490 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  1.760 1.635 3.620 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.465 0.780 5.760 0.890 ;
        RECT  5.370 0.555 5.465 1.525 ;
        RECT  5.355 0.555 5.370 0.665 ;
        RECT  5.305 1.315 5.370 1.525 ;
        RECT  5.245 0.285 5.355 0.665 ;
        RECT  5.190 0.780 5.280 0.890 ;
        RECT  5.000 0.555 5.245 0.665 ;
        RECT  5.100 0.780 5.190 1.305 ;
        RECT  4.170 1.215 5.100 1.305 ;
        RECT  4.890 0.555 5.000 0.920 ;
        RECT  4.500 1.015 4.965 1.125 ;
        RECT  4.500 0.275 4.655 0.405 ;
        RECT  4.410 0.275 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  3.105 0.275 4.320 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  3.335 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.045 1.015 3.575 1.125 ;
        RECT  3.230 0.495 3.340 0.905 ;
        RECT  3.245 1.215 3.335 1.525 ;
        RECT  2.635 1.425 3.245 1.525 ;
        RECT  2.700 0.495 3.230 0.605 ;
        RECT  2.745 0.275 3.105 0.365 ;
        RECT  2.935 0.900 3.045 1.125 ;
        RECT  2.590 0.495 2.700 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.275 1.295 2.445 1.445 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.065 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  1.460 1.295 2.275 1.385 ;
        RECT  1.960 0.800 2.135 0.910 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSNQD1

MACRO SDFSNQD2
    CLASS CORE ;
    FOREIGN SDFSNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0790 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.630 0.510 4.750 0.925 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 0.285 5.950 1.490 ;
        RECT  5.765 0.285 5.850 0.665 ;
        RECT  5.765 1.050 5.850 1.490 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.080 -0.165 6.200 0.165 ;
        RECT  4.970 -0.165 5.080 0.465 ;
        RECT  0.520 -0.165 4.970 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.090 1.635 6.200 1.965 ;
        RECT  4.980 1.455 5.090 1.965 ;
        RECT  4.620 1.635 4.980 1.965 ;
        RECT  4.450 1.395 4.620 1.965 ;
        RECT  3.705 1.635 4.450 1.965 ;
        RECT  3.595 1.395 3.705 1.965 ;
        RECT  1.760 1.635 3.595 1.965 ;
        RECT  1.570 1.495 1.760 1.965 ;
        RECT  0.470 1.635 1.570 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.500 0.780 5.760 0.890 ;
        RECT  5.410 0.555 5.500 1.150 ;
        RECT  5.345 0.555 5.410 0.665 ;
        RECT  5.375 1.050 5.410 1.150 ;
        RECT  5.265 1.050 5.375 1.460 ;
        RECT  5.235 0.285 5.345 0.665 ;
        RECT  5.175 0.780 5.320 0.890 ;
        RECT  4.985 0.555 5.235 0.665 ;
        RECT  5.085 0.780 5.175 1.305 ;
        RECT  4.140 1.215 5.085 1.305 ;
        RECT  4.875 0.555 4.985 0.920 ;
        RECT  4.500 1.015 4.925 1.125 ;
        RECT  4.500 0.310 4.665 0.420 ;
        RECT  4.410 0.310 4.500 1.125 ;
        RECT  4.050 0.545 4.410 0.655 ;
        RECT  4.245 1.015 4.410 1.125 ;
        RECT  2.745 0.275 4.305 0.375 ;
        RECT  4.040 0.835 4.140 1.305 ;
        RECT  3.930 0.835 4.040 0.925 ;
        RECT  3.820 0.495 3.930 0.925 ;
        RECT  3.825 1.215 3.930 1.525 ;
        RECT  3.670 1.015 3.910 1.125 ;
        RECT  3.320 1.215 3.825 1.305 ;
        RECT  3.560 0.495 3.670 1.125 ;
        RECT  3.040 1.015 3.560 1.125 ;
        RECT  3.215 0.495 3.325 0.905 ;
        RECT  3.230 1.215 3.320 1.525 ;
        RECT  2.630 1.425 3.230 1.525 ;
        RECT  2.695 0.495 3.215 0.605 ;
        RECT  2.930 0.900 3.040 1.125 ;
        RECT  2.585 0.495 2.695 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.280 1.295 2.430 1.490 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.060 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  1.460 1.295 2.280 1.385 ;
        RECT  1.960 0.780 2.135 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.295 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSNQD2

MACRO SDFSNQD4
    CLASS CORE ;
    FOREIGN SDFSNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.815 0.600 1.090 ;
        RECT  0.445 0.700 0.555 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0644 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.700 0.175 1.090 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0790 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.630 0.510 4.760 0.925 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.325 6.475 0.635 ;
        RECT  6.250 1.100 6.475 1.410 ;
        RECT  5.950 0.325 6.250 1.410 ;
        RECT  5.805 0.325 5.950 0.640 ;
        RECT  5.805 1.100 5.950 1.410 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.710 1.355 1.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.705 -0.165 6.800 0.165 ;
        RECT  6.595 -0.165 6.705 0.685 ;
        RECT  5.685 -0.165 6.595 0.165 ;
        RECT  5.575 -0.165 5.685 0.465 ;
        RECT  5.130 -0.165 5.575 0.165 ;
        RECT  5.020 -0.165 5.130 0.465 ;
        RECT  0.520 -0.165 5.020 0.165 ;
        RECT  0.310 -0.165 0.520 0.400 ;
        RECT  0.000 -0.165 0.310 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.705 1.635 6.800 1.965 ;
        RECT  6.595 1.050 6.705 1.965 ;
        RECT  5.685 1.635 6.595 1.965 ;
        RECT  5.575 1.250 5.685 1.965 ;
        RECT  4.665 1.635 5.575 1.965 ;
        RECT  4.495 1.395 4.665 1.965 ;
        RECT  3.730 1.635 4.495 1.965 ;
        RECT  3.620 1.395 3.730 1.965 ;
        RECT  0.470 1.635 3.620 1.965 ;
        RECT  0.360 1.380 0.470 1.965 ;
        RECT  0.000 1.635 0.360 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.350 0.325 6.475 0.635 ;
        RECT  6.350 1.100 6.475 1.410 ;
        RECT  5.805 0.325 5.850 0.640 ;
        RECT  5.805 1.100 5.850 1.410 ;
        RECT  5.495 0.785 5.840 0.890 ;
        RECT  5.425 0.555 5.495 1.150 ;
        RECT  5.405 0.555 5.425 1.460 ;
        RECT  5.395 0.555 5.405 0.665 ;
        RECT  5.315 1.050 5.405 1.460 ;
        RECT  5.285 0.285 5.395 0.665 ;
        RECT  5.225 0.780 5.315 0.890 ;
        RECT  5.035 0.555 5.285 0.665 ;
        RECT  5.135 0.780 5.225 1.305 ;
        RECT  4.170 1.215 5.135 1.305 ;
        RECT  4.925 0.555 5.035 0.920 ;
        RECT  4.500 1.015 4.975 1.125 ;
        RECT  4.500 0.310 4.705 0.420 ;
        RECT  4.410 0.310 4.500 1.125 ;
        RECT  4.065 0.545 4.410 0.655 ;
        RECT  4.275 1.015 4.410 1.125 ;
        RECT  3.105 0.275 4.320 0.375 ;
        RECT  4.070 0.835 4.170 1.305 ;
        RECT  3.945 0.835 4.070 0.925 ;
        RECT  3.855 1.215 3.960 1.525 ;
        RECT  3.835 0.495 3.945 0.925 ;
        RECT  3.685 1.015 3.940 1.125 ;
        RECT  3.335 1.215 3.855 1.305 ;
        RECT  3.575 0.495 3.685 1.125 ;
        RECT  3.045 1.015 3.575 1.125 ;
        RECT  3.230 0.495 3.340 0.905 ;
        RECT  3.245 1.215 3.335 1.525 ;
        RECT  2.635 1.425 3.245 1.525 ;
        RECT  2.700 0.495 3.230 0.605 ;
        RECT  2.745 0.275 3.105 0.365 ;
        RECT  2.935 0.900 3.045 1.125 ;
        RECT  2.590 0.495 2.700 1.315 ;
        RECT  2.335 0.295 2.550 0.405 ;
        RECT  1.460 1.335 2.465 1.445 ;
        RECT  2.340 0.545 2.450 1.145 ;
        RECT  2.110 0.545 2.340 0.655 ;
        RECT  2.060 1.035 2.340 1.145 ;
        RECT  0.865 0.305 2.335 0.405 ;
        RECT  1.960 0.780 2.135 0.890 ;
        RECT  1.860 0.510 1.960 1.195 ;
        RECT  1.615 0.510 1.860 0.620 ;
        RECT  1.555 1.085 1.860 1.195 ;
        RECT  1.360 1.335 1.460 1.525 ;
        RECT  0.945 1.435 1.360 1.525 ;
        RECT  1.140 0.500 1.325 0.600 ;
        RECT  1.140 1.215 1.250 1.325 ;
        RECT  1.050 0.500 1.140 1.325 ;
        RECT  0.835 1.135 0.945 1.525 ;
        RECT  0.750 0.595 0.850 0.915 ;
        RECT  0.740 0.490 0.750 0.915 ;
        RECT  0.660 0.490 0.740 0.705 ;
        RECT  0.355 0.490 0.660 0.590 ;
        RECT  0.265 0.490 0.355 1.290 ;
        RECT  0.185 0.490 0.265 0.590 ;
        RECT  0.185 1.200 0.265 1.290 ;
        RECT  0.075 0.385 0.185 0.590 ;
        RECT  0.075 1.200 0.185 1.450 ;
    END
END SDFSNQD4

MACRO SDFXD0
    CLASS CORE ;
    FOREIGN SDFXD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0183 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0521 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 0.890 ;
        RECT  0.430 0.670 0.450 0.890 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0449 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.000 2.950 1.290 ;
        RECT  2.780 1.000 2.850 1.090 ;
        RECT  2.650 0.910 2.780 1.090 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.475 7.150 1.290 ;
        RECT  7.020 0.475 7.050 0.665 ;
        RECT  7.015 1.020 7.050 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.630 6.750 1.120 ;
        RECT  6.625 0.630 6.650 0.730 ;
        RECT  6.625 1.020 6.650 1.120 ;
        RECT  6.525 0.475 6.625 0.730 ;
        RECT  6.525 1.020 6.625 1.230 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0227 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.890 2.350 1.090 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0321 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.890 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.850 4.350 1.290 ;
        RECT  4.160 0.850 4.250 1.020 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.790 -0.165 7.200 0.165 ;
        RECT  4.680 -0.165 4.790 0.420 ;
        RECT  0.185 -0.165 4.680 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.840 1.635 7.200 1.965 ;
        RECT  6.730 1.455 6.840 1.965 ;
        RECT  3.880 1.635 6.730 1.965 ;
        RECT  3.770 1.335 3.880 1.965 ;
        RECT  0.000 1.635 3.770 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.930 0.735 6.960 0.905 ;
        RECT  6.840 0.275 6.930 0.905 ;
        RECT  6.365 0.275 6.840 0.365 ;
        RECT  6.365 0.615 6.435 1.370 ;
        RECT  6.345 0.275 6.365 1.370 ;
        RECT  6.255 0.275 6.345 0.725 ;
        RECT  6.225 1.260 6.345 1.370 ;
        RECT  5.870 0.615 6.255 0.725 ;
        RECT  6.005 0.945 6.255 1.055 ;
        RECT  5.915 0.825 6.005 1.345 ;
        RECT  5.780 0.825 5.915 0.915 ;
        RECT  5.520 1.235 5.915 1.345 ;
        RECT  5.690 0.305 5.780 0.915 ;
        RECT  5.430 1.005 5.775 1.105 ;
        RECT  5.510 0.305 5.690 0.415 ;
        RECT  5.430 0.565 5.595 0.675 ;
        RECT  5.325 1.435 5.535 1.545 ;
        RECT  5.340 0.565 5.430 1.320 ;
        RECT  4.740 0.580 5.340 0.690 ;
        RECT  4.725 1.210 5.340 1.320 ;
        RECT  5.030 1.435 5.325 1.525 ;
        RECT  5.125 0.830 5.235 1.120 ;
        RECT  4.635 1.030 5.125 1.120 ;
        RECT  4.815 1.435 5.030 1.545 ;
        RECT  4.125 1.435 4.815 1.525 ;
        RECT  4.620 1.030 4.635 1.305 ;
        RECT  4.510 0.615 4.620 1.305 ;
        RECT  4.440 0.275 4.550 0.525 ;
        RECT  4.350 0.615 4.510 0.715 ;
        RECT  3.385 0.275 4.440 0.365 ;
        RECT  4.260 0.455 4.350 0.715 ;
        RECT  3.730 0.455 4.260 0.545 ;
        RECT  4.070 0.645 4.170 0.755 ;
        RECT  4.070 1.300 4.125 1.525 ;
        RECT  3.980 0.645 4.070 1.525 ;
        RECT  3.350 1.055 3.980 1.165 ;
        RECT  3.620 0.455 3.730 0.935 ;
        RECT  3.275 0.275 3.385 0.535 ;
        RECT  3.265 1.255 3.375 1.525 ;
        RECT  3.260 0.625 3.350 1.165 ;
        RECT  3.050 0.445 3.275 0.535 ;
        RECT  3.150 1.255 3.265 1.345 ;
        RECT  3.160 0.625 3.260 0.725 ;
        RECT  3.060 0.820 3.150 1.345 ;
        RECT  1.895 1.435 3.140 1.525 ;
        RECT  2.870 0.265 3.130 0.355 ;
        RECT  3.050 0.820 3.060 0.910 ;
        RECT  2.960 0.445 3.050 0.910 ;
        RECT  2.760 0.265 2.870 0.365 ;
        RECT  0.665 0.275 2.760 0.365 ;
        RECT  2.560 1.215 2.675 1.325 ;
        RECT  2.560 0.465 2.625 0.800 ;
        RECT  2.515 0.465 2.560 1.325 ;
        RECT  2.470 0.700 2.515 1.325 ;
        RECT  1.945 0.700 2.470 0.800 ;
        RECT  1.230 0.495 2.395 0.585 ;
        RECT  1.215 1.205 2.380 1.315 ;
        RECT  1.855 0.700 1.945 1.095 ;
        RECT  1.685 1.405 1.895 1.525 ;
        RECT  1.320 1.000 1.855 1.095 ;
        RECT  0.625 1.435 1.685 1.525 ;
        RECT  0.895 0.725 1.290 0.835 ;
        RECT  0.875 0.470 0.895 1.100 ;
        RECT  0.785 0.470 0.875 1.345 ;
        RECT  0.765 0.990 0.785 1.345 ;
        RECT  0.390 0.990 0.765 1.100 ;
        RECT  0.475 0.275 0.665 0.405 ;
        RECT  0.515 1.255 0.625 1.525 ;
    END
END SDFXD0

MACRO SDFXD1
    CLASS CORE ;
    FOREIGN SDFXD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0583 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 0.890 ;
        RECT  0.430 0.670 0.450 0.890 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0650 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.000 2.950 1.290 ;
        RECT  2.780 1.000 2.850 1.090 ;
        RECT  2.650 0.910 2.780 1.090 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.275 7.150 1.490 ;
        RECT  7.020 0.275 7.050 0.665 ;
        RECT  7.015 1.050 7.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.630 6.750 1.120 ;
        RECT  6.625 0.630 6.650 0.730 ;
        RECT  6.625 1.020 6.650 1.120 ;
        RECT  6.525 0.475 6.625 0.730 ;
        RECT  6.525 1.020 6.625 1.460 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.890 2.350 1.090 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0322 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.890 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.850 4.350 1.290 ;
        RECT  4.160 0.850 4.250 1.020 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.790 -0.165 7.200 0.165 ;
        RECT  4.680 -0.165 4.790 0.420 ;
        RECT  0.185 -0.165 4.680 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.880 1.635 7.200 1.965 ;
        RECT  3.770 1.335 3.880 1.965 ;
        RECT  0.185 1.635 3.770 1.965 ;
        RECT  0.075 1.280 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.930 0.735 6.960 0.905 ;
        RECT  6.840 0.275 6.930 0.905 ;
        RECT  6.365 0.275 6.840 0.365 ;
        RECT  6.365 0.615 6.435 1.410 ;
        RECT  6.345 0.275 6.365 1.410 ;
        RECT  6.255 0.275 6.345 0.725 ;
        RECT  6.235 1.300 6.345 1.410 ;
        RECT  5.870 0.615 6.255 0.725 ;
        RECT  6.005 0.945 6.255 1.055 ;
        RECT  5.915 0.825 6.005 1.345 ;
        RECT  5.780 0.825 5.915 0.915 ;
        RECT  5.520 1.235 5.915 1.345 ;
        RECT  5.690 0.305 5.780 0.915 ;
        RECT  5.430 1.005 5.775 1.105 ;
        RECT  5.510 0.305 5.690 0.415 ;
        RECT  5.430 0.565 5.595 0.675 ;
        RECT  5.325 1.435 5.535 1.545 ;
        RECT  5.340 0.565 5.430 1.320 ;
        RECT  4.740 0.580 5.340 0.690 ;
        RECT  4.725 1.210 5.340 1.320 ;
        RECT  5.030 1.435 5.325 1.525 ;
        RECT  5.125 0.830 5.235 1.120 ;
        RECT  4.635 1.030 5.125 1.120 ;
        RECT  4.815 1.435 5.030 1.545 ;
        RECT  4.125 1.435 4.815 1.525 ;
        RECT  4.620 1.030 4.635 1.305 ;
        RECT  4.510 0.615 4.620 1.305 ;
        RECT  4.440 0.275 4.550 0.525 ;
        RECT  4.350 0.615 4.510 0.715 ;
        RECT  3.385 0.275 4.440 0.365 ;
        RECT  4.260 0.455 4.350 0.715 ;
        RECT  3.730 0.455 4.260 0.545 ;
        RECT  4.070 0.635 4.170 0.745 ;
        RECT  4.070 1.120 4.125 1.525 ;
        RECT  3.980 0.635 4.070 1.525 ;
        RECT  3.350 1.055 3.980 1.165 ;
        RECT  3.620 0.455 3.730 0.935 ;
        RECT  3.275 0.275 3.385 0.535 ;
        RECT  3.265 1.255 3.375 1.525 ;
        RECT  3.260 0.625 3.350 1.165 ;
        RECT  3.050 0.445 3.275 0.535 ;
        RECT  3.150 1.255 3.265 1.345 ;
        RECT  3.160 0.625 3.260 0.725 ;
        RECT  3.060 0.820 3.150 1.345 ;
        RECT  1.915 1.435 3.140 1.525 ;
        RECT  2.870 0.265 3.130 0.355 ;
        RECT  3.050 0.820 3.060 0.910 ;
        RECT  2.960 0.445 3.050 0.910 ;
        RECT  2.760 0.265 2.870 0.365 ;
        RECT  0.665 0.275 2.760 0.365 ;
        RECT  2.560 1.215 2.675 1.325 ;
        RECT  2.560 0.455 2.625 0.800 ;
        RECT  2.515 0.455 2.560 1.325 ;
        RECT  2.470 0.700 2.515 1.325 ;
        RECT  1.945 0.700 2.470 0.800 ;
        RECT  1.230 0.495 2.395 0.585 ;
        RECT  1.235 1.205 2.380 1.315 ;
        RECT  1.855 0.700 1.945 1.095 ;
        RECT  1.705 1.405 1.915 1.525 ;
        RECT  1.340 1.000 1.855 1.095 ;
        RECT  0.635 1.435 1.705 1.525 ;
        RECT  0.900 0.725 1.290 0.835 ;
        RECT  0.785 0.470 0.900 1.345 ;
        RECT  0.400 0.990 0.785 1.100 ;
        RECT  0.475 0.275 0.665 0.405 ;
        RECT  0.525 1.275 0.635 1.525 ;
    END
END SDFXD1

MACRO SDFXD2
    CLASS CORE ;
    FOREIGN SDFXD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0583 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 0.890 ;
        RECT  0.430 0.670 0.450 0.890 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0650 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.000 2.950 1.290 ;
        RECT  2.780 1.000 2.850 1.090 ;
        RECT  2.650 0.910 2.780 1.090 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.565 7.550 1.150 ;
        RECT  7.445 0.565 7.450 0.665 ;
        RECT  7.445 1.050 7.450 1.150 ;
        RECT  7.335 0.275 7.445 0.665 ;
        RECT  7.335 1.050 7.445 1.460 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.475 6.950 1.490 ;
        RECT  6.815 0.475 6.850 0.685 ;
        RECT  6.815 1.020 6.850 1.490 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.890 2.350 1.090 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0322 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.890 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.850 4.350 1.290 ;
        RECT  4.160 0.850 4.250 1.020 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 -0.165 7.800 0.165 ;
        RECT  7.595 -0.165 7.705 0.485 ;
        RECT  6.135 -0.165 7.595 0.165 ;
        RECT  6.025 -0.165 6.135 0.465 ;
        RECT  4.790 -0.165 6.025 0.165 ;
        RECT  4.680 -0.165 4.790 0.420 ;
        RECT  0.185 -0.165 4.680 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 1.635 7.800 1.965 ;
        RECT  7.595 1.250 7.705 1.965 ;
        RECT  7.185 1.635 7.595 1.965 ;
        RECT  7.075 1.050 7.185 1.965 ;
        RECT  6.665 1.635 7.075 1.965 ;
        RECT  6.555 1.050 6.665 1.965 ;
        RECT  3.880 1.635 6.555 1.965 ;
        RECT  3.770 1.335 3.880 1.965 ;
        RECT  0.185 1.635 3.770 1.965 ;
        RECT  0.075 1.275 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.180 0.765 7.360 0.875 ;
        RECT  7.090 0.275 7.180 0.875 ;
        RECT  6.395 0.275 7.090 0.365 ;
        RECT  6.395 0.615 6.465 1.410 ;
        RECT  6.375 0.275 6.395 1.410 ;
        RECT  6.285 0.275 6.375 0.725 ;
        RECT  6.225 1.300 6.375 1.410 ;
        RECT  5.870 0.615 6.285 0.725 ;
        RECT  6.005 0.945 6.285 1.055 ;
        RECT  5.915 0.825 6.005 1.345 ;
        RECT  5.780 0.825 5.915 0.915 ;
        RECT  5.520 1.235 5.915 1.345 ;
        RECT  5.690 0.305 5.780 0.915 ;
        RECT  5.430 1.005 5.775 1.105 ;
        RECT  5.510 0.305 5.690 0.415 ;
        RECT  5.430 0.565 5.595 0.675 ;
        RECT  5.325 1.435 5.535 1.545 ;
        RECT  5.340 0.565 5.430 1.320 ;
        RECT  4.740 0.580 5.340 0.690 ;
        RECT  4.725 1.210 5.340 1.320 ;
        RECT  5.030 1.435 5.325 1.525 ;
        RECT  5.125 0.830 5.235 1.120 ;
        RECT  4.635 1.030 5.125 1.120 ;
        RECT  4.815 1.435 5.030 1.545 ;
        RECT  4.125 1.435 4.815 1.525 ;
        RECT  4.620 1.030 4.635 1.305 ;
        RECT  4.510 0.615 4.620 1.305 ;
        RECT  4.440 0.275 4.550 0.525 ;
        RECT  4.350 0.615 4.510 0.715 ;
        RECT  3.385 0.275 4.440 0.365 ;
        RECT  4.260 0.455 4.350 0.715 ;
        RECT  3.730 0.455 4.260 0.545 ;
        RECT  4.070 0.635 4.170 0.745 ;
        RECT  4.070 1.120 4.125 1.525 ;
        RECT  3.980 0.635 4.070 1.525 ;
        RECT  3.350 1.055 3.980 1.165 ;
        RECT  3.620 0.455 3.730 0.935 ;
        RECT  3.275 0.275 3.385 0.535 ;
        RECT  3.265 1.255 3.375 1.525 ;
        RECT  3.260 0.625 3.350 1.165 ;
        RECT  3.050 0.445 3.275 0.535 ;
        RECT  3.150 1.255 3.265 1.345 ;
        RECT  3.160 0.625 3.260 0.725 ;
        RECT  3.060 0.820 3.150 1.345 ;
        RECT  1.915 1.435 3.140 1.525 ;
        RECT  2.870 0.265 3.130 0.355 ;
        RECT  3.050 0.820 3.060 0.910 ;
        RECT  2.960 0.445 3.050 0.910 ;
        RECT  2.760 0.265 2.870 0.365 ;
        RECT  0.665 0.275 2.760 0.365 ;
        RECT  2.560 1.215 2.675 1.325 ;
        RECT  2.560 0.455 2.625 0.800 ;
        RECT  2.515 0.455 2.560 1.325 ;
        RECT  2.470 0.700 2.515 1.325 ;
        RECT  1.945 0.700 2.470 0.800 ;
        RECT  1.230 0.495 2.395 0.585 ;
        RECT  1.235 1.205 2.380 1.315 ;
        RECT  1.855 0.700 1.945 1.095 ;
        RECT  1.705 1.405 1.915 1.525 ;
        RECT  1.340 1.000 1.855 1.095 ;
        RECT  0.635 1.435 1.705 1.525 ;
        RECT  0.900 0.725 1.290 0.835 ;
        RECT  0.785 0.470 0.900 1.345 ;
        RECT  0.400 0.990 0.785 1.100 ;
        RECT  0.475 0.275 0.665 0.405 ;
        RECT  0.525 1.270 0.635 1.525 ;
    END
END SDFXD2

MACRO SDFXD4
    CLASS CORE ;
    FOREIGN SDFXD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0583 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 0.890 ;
        RECT  0.430 0.670 0.450 0.890 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0650 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.000 2.950 1.290 ;
        RECT  2.780 1.000 2.850 1.090 ;
        RECT  2.650 0.910 2.780 1.090 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.850 0.325 9.075 0.635 ;
        RECT  8.850 1.100 9.075 1.410 ;
        RECT  8.550 0.325 8.850 1.410 ;
        RECT  8.405 0.325 8.550 0.635 ;
        RECT  8.405 1.100 8.550 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 0.325 8.055 0.635 ;
        RECT  7.850 1.110 8.050 1.290 ;
        RECT  7.550 0.325 7.850 1.290 ;
        RECT  7.385 0.325 7.550 0.635 ;
        RECT  7.370 1.110 7.550 1.290 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.890 2.350 1.090 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0322 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.890 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0445 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.910 4.150 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.305 -0.165 9.400 0.165 ;
        RECT  9.195 -0.165 9.305 0.685 ;
        RECT  8.285 -0.165 9.195 0.165 ;
        RECT  8.175 -0.165 8.285 0.665 ;
        RECT  6.810 -0.165 8.175 0.165 ;
        RECT  6.640 -0.165 6.810 0.415 ;
        RECT  5.770 -0.165 6.640 0.165 ;
        RECT  5.600 -0.165 5.770 0.405 ;
        RECT  4.715 -0.165 5.600 0.165 ;
        RECT  4.605 -0.165 4.715 0.725 ;
        RECT  3.940 -0.165 4.605 0.165 ;
        RECT  3.770 -0.165 3.940 0.355 ;
        RECT  0.185 -0.165 3.770 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.305 1.635 9.400 1.965 ;
        RECT  9.195 1.050 9.305 1.965 ;
        RECT  5.880 1.635 9.195 1.965 ;
        RECT  5.790 1.135 5.880 1.965 ;
        RECT  5.625 1.135 5.790 1.245 ;
        RECT  0.185 1.635 5.790 1.965 ;
        RECT  0.075 1.275 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.950 0.325 9.075 0.635 ;
        RECT  8.950 1.100 9.075 1.410 ;
        RECT  8.405 0.325 8.450 0.635 ;
        RECT  8.405 1.100 8.450 1.410 ;
        RECT  7.950 0.325 8.055 0.635 ;
        RECT  7.950 1.110 8.050 1.290 ;
        RECT  7.385 0.325 7.450 0.635 ;
        RECT  7.370 1.110 7.450 1.290 ;
        RECT  8.295 0.780 8.440 0.890 ;
        RECT  8.185 0.780 8.295 1.505 ;
        RECT  7.195 1.395 8.185 1.505 ;
        RECT  7.105 0.585 7.195 1.505 ;
        RECT  7.055 0.585 7.105 0.675 ;
        RECT  6.940 1.105 7.105 1.505 ;
        RECT  6.935 0.275 7.055 0.675 ;
        RECT  6.715 0.780 7.005 0.890 ;
        RECT  6.645 0.585 6.935 0.675 ;
        RECT  6.610 0.780 6.715 1.500 ;
        RECT  6.535 0.505 6.645 0.675 ;
        RECT  6.420 0.780 6.610 0.890 ;
        RECT  6.060 1.390 6.610 1.500 ;
        RECT  6.340 1.060 6.450 1.280 ;
        RECT  6.330 0.305 6.420 0.890 ;
        RECT  6.240 1.060 6.340 1.160 ;
        RECT  5.965 0.305 6.330 0.415 ;
        RECT  6.190 0.735 6.240 1.160 ;
        RECT  6.150 0.560 6.190 1.160 ;
        RECT  6.080 0.560 6.150 0.845 ;
        RECT  4.975 0.735 6.080 0.845 ;
        RECT  5.970 0.955 6.060 1.500 ;
        RECT  5.480 0.955 5.970 1.045 ;
        RECT  5.875 0.305 5.965 0.605 ;
        RECT  5.235 0.495 5.875 0.605 ;
        RECT  5.480 1.345 5.700 1.515 ;
        RECT  5.370 0.955 5.480 1.165 ;
        RECT  5.370 1.255 5.480 1.515 ;
        RECT  5.185 1.055 5.370 1.165 ;
        RECT  4.705 1.255 5.370 1.345 ;
        RECT  5.065 1.435 5.240 1.545 ;
        RECT  5.125 0.335 5.235 0.605 ;
        RECT  4.975 1.055 5.095 1.165 ;
        RECT  4.375 1.435 5.065 1.525 ;
        RECT  4.865 0.490 4.975 1.165 ;
        RECT  4.580 1.175 4.705 1.345 ;
        RECT  4.480 1.175 4.580 1.285 ;
        RECT  4.165 0.305 4.480 0.415 ;
        RECT  4.390 0.515 4.480 1.285 ;
        RECT  4.345 0.515 4.390 0.725 ;
        RECT  3.760 1.180 4.390 1.285 ;
        RECT  4.245 1.385 4.375 1.525 ;
        RECT  3.560 1.385 4.245 1.495 ;
        RECT  3.560 0.625 4.225 0.735 ;
        RECT  4.075 0.305 4.165 0.535 ;
        RECT  3.445 0.445 4.075 0.535 ;
        RECT  3.670 0.915 3.760 1.285 ;
        RECT  3.470 0.625 3.560 1.495 ;
        RECT  3.175 0.625 3.470 0.735 ;
        RECT  3.420 1.075 3.470 1.245 ;
        RECT  3.315 0.275 3.445 0.535 ;
        RECT  3.310 1.355 3.365 1.525 ;
        RECT  3.085 0.445 3.315 0.535 ;
        RECT  3.210 0.825 3.310 1.525 ;
        RECT  3.085 0.825 3.210 0.915 ;
        RECT  2.865 0.265 3.130 0.355 ;
        RECT  3.005 1.365 3.115 1.545 ;
        RECT  2.995 0.445 3.085 0.915 ;
        RECT  1.915 1.435 3.005 1.525 ;
        RECT  2.760 0.265 2.865 0.365 ;
        RECT  0.665 0.275 2.760 0.365 ;
        RECT  2.560 1.215 2.675 1.325 ;
        RECT  2.560 0.455 2.625 0.800 ;
        RECT  2.515 0.455 2.560 1.325 ;
        RECT  2.470 0.700 2.515 1.325 ;
        RECT  1.945 0.700 2.470 0.800 ;
        RECT  1.230 0.495 2.395 0.585 ;
        RECT  1.235 1.205 2.380 1.315 ;
        RECT  1.855 0.700 1.945 1.095 ;
        RECT  1.705 1.405 1.915 1.525 ;
        RECT  1.340 1.000 1.855 1.095 ;
        RECT  0.635 1.435 1.705 1.525 ;
        RECT  0.900 0.725 1.290 0.835 ;
        RECT  0.785 0.470 0.900 1.345 ;
        RECT  0.400 0.990 0.785 1.100 ;
        RECT  0.475 0.275 0.665 0.405 ;
        RECT  0.525 1.275 0.635 1.525 ;
    END
END SDFXD4

MACRO SDFXQD0
    CLASS CORE ;
    FOREIGN SDFXQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.710 3.150 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0483 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.710 1.750 1.090 ;
        RECT  1.530 0.845 1.650 1.015 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0471 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END SA
    PIN Q
        ANTENNAGATEAREA 0.0180 ;
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.430 6.150 1.490 ;
        RECT  6.015 0.430 6.050 0.720 ;
        RECT  6.015 1.280 6.050 1.490 ;
        RECT  5.775 0.610 6.015 0.720 ;
        RECT  5.675 0.610 5.775 0.875 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0261 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.510 1.010 0.700 ;
        RECT  0.850 0.510 0.950 0.890 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0261 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.750 0.700 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.710 3.460 0.890 ;
        RECT  3.250 0.710 3.350 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.165 6.200 0.165 ;
        RECT  1.805 -0.165 1.910 0.425 ;
        RECT  0.000 -0.165 1.805 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.635 6.200 1.965 ;
        RECT  4.735 1.350 4.845 1.965 ;
        RECT  0.525 1.635 4.735 1.965 ;
        RECT  0.435 1.200 0.525 1.965 ;
        RECT  0.300 1.200 0.435 1.310 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.850 0.995 5.960 1.190 ;
        RECT  5.805 1.100 5.850 1.190 ;
        RECT  5.705 1.100 5.805 1.495 ;
        RECT  5.360 1.385 5.705 1.495 ;
        RECT  5.495 0.275 5.585 1.295 ;
        RECT  5.340 0.275 5.495 0.365 ;
        RECT  5.450 1.085 5.495 1.295 ;
        RECT  5.360 0.455 5.405 0.665 ;
        RECT  5.270 0.455 5.360 1.495 ;
        RECT  5.170 0.255 5.340 0.365 ;
        RECT  5.250 1.385 5.270 1.495 ;
        RECT  5.090 0.455 5.180 1.245 ;
        RECT  4.590 0.275 5.170 0.365 ;
        RECT  5.040 0.455 5.090 0.645 ;
        RECT  4.770 1.135 5.090 1.245 ;
        RECT  4.950 0.735 5.000 0.905 ;
        RECT  4.860 0.465 4.950 0.905 ;
        RECT  4.500 0.465 4.860 0.555 ;
        RECT  4.670 0.735 4.770 1.245 ;
        RECT  4.420 0.255 4.590 0.365 ;
        RECT  4.410 0.465 4.500 1.085 ;
        RECT  4.300 0.465 4.410 0.565 ;
        RECT  4.360 0.985 4.410 1.085 ;
        RECT  4.250 0.985 4.360 1.265 ;
        RECT  4.050 0.765 4.205 0.875 ;
        RECT  3.990 0.255 4.160 0.365 ;
        RECT  3.960 1.235 4.130 1.525 ;
        RECT  3.955 0.505 4.050 1.135 ;
        RECT  2.395 0.275 3.990 0.365 ;
        RECT  2.390 1.435 3.960 1.525 ;
        RECT  3.775 0.505 3.955 0.615 ;
        RECT  3.745 1.025 3.955 1.135 ;
        RECT  3.655 0.770 3.830 0.880 ;
        RECT  3.565 0.505 3.655 1.290 ;
        RECT  3.245 0.505 3.565 0.615 ;
        RECT  3.225 1.180 3.565 1.290 ;
        RECT  2.730 0.485 3.155 0.595 ;
        RECT  3.005 1.000 3.115 1.315 ;
        RECT  2.730 1.000 3.005 1.110 ;
        RECT  2.620 0.485 2.730 1.110 ;
        RECT  2.380 0.730 2.490 1.085 ;
        RECT  2.285 0.275 2.395 0.625 ;
        RECT  2.280 1.215 2.390 1.525 ;
        RECT  2.010 0.730 2.380 0.820 ;
        RECT  2.190 0.945 2.290 1.055 ;
        RECT  2.100 0.945 2.190 1.525 ;
        RECT  1.440 1.435 2.100 1.525 ;
        RECT  1.900 0.515 2.010 1.325 ;
        RECT  1.645 0.515 1.900 0.605 ;
        RECT  1.555 1.215 1.900 1.325 ;
        RECT  1.535 0.265 1.645 0.605 ;
        RECT  1.350 0.310 1.440 1.525 ;
        RECT  0.775 0.310 1.350 0.420 ;
        RECT  0.765 1.210 1.350 1.300 ;
        RECT  1.150 0.515 1.260 1.090 ;
        RECT  0.750 1.000 1.150 1.090 ;
        RECT  0.660 0.885 0.750 1.090 ;
        RECT  0.360 0.885 0.660 0.995 ;
        RECT  0.270 0.305 0.360 1.090 ;
        RECT  0.045 0.305 0.270 0.415 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.320 ;
    END
END SDFXQD0

MACRO SDFXQD1
    CLASS CORE ;
    FOREIGN SDFXQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0583 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 0.890 ;
        RECT  0.430 0.670 0.450 0.890 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0650 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.000 2.950 1.290 ;
        RECT  2.780 1.000 2.850 1.090 ;
        RECT  2.650 0.910 2.780 1.090 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.275 6.950 1.490 ;
        RECT  6.775 0.275 6.850 0.685 ;
        RECT  6.775 1.050 6.850 1.490 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.890 2.350 1.090 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0322 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.890 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.850 4.350 1.290 ;
        RECT  4.160 0.850 4.250 1.020 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.625 -0.165 7.000 0.165 ;
        RECT  6.515 -0.165 6.625 0.505 ;
        RECT  4.790 -0.165 6.515 0.165 ;
        RECT  4.680 -0.165 4.790 0.420 ;
        RECT  0.185 -0.165 4.680 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.625 1.635 7.000 1.965 ;
        RECT  6.515 1.335 6.625 1.965 ;
        RECT  3.880 1.635 6.515 1.965 ;
        RECT  3.770 1.335 3.880 1.965 ;
        RECT  0.185 1.635 3.770 1.965 ;
        RECT  0.075 1.275 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.575 0.615 6.665 1.245 ;
        RECT  6.365 0.615 6.575 0.725 ;
        RECT  6.375 1.155 6.575 1.245 ;
        RECT  6.265 1.155 6.375 1.375 ;
        RECT  6.255 0.255 6.365 0.725 ;
        RECT  5.870 0.615 6.255 0.725 ;
        RECT  6.005 0.945 6.255 1.055 ;
        RECT  5.915 0.825 6.005 1.345 ;
        RECT  5.780 0.825 5.915 0.915 ;
        RECT  5.520 1.235 5.915 1.345 ;
        RECT  5.690 0.305 5.780 0.915 ;
        RECT  5.430 1.005 5.775 1.105 ;
        RECT  5.510 0.305 5.690 0.415 ;
        RECT  5.430 0.565 5.595 0.675 ;
        RECT  5.325 1.435 5.535 1.545 ;
        RECT  5.340 0.565 5.430 1.320 ;
        RECT  4.740 0.580 5.340 0.690 ;
        RECT  4.725 1.210 5.340 1.320 ;
        RECT  5.030 1.435 5.325 1.525 ;
        RECT  5.125 0.830 5.235 1.120 ;
        RECT  4.635 1.030 5.125 1.120 ;
        RECT  4.815 1.435 5.030 1.545 ;
        RECT  4.125 1.435 4.815 1.525 ;
        RECT  4.620 1.030 4.635 1.305 ;
        RECT  4.510 0.615 4.620 1.305 ;
        RECT  4.440 0.275 4.550 0.525 ;
        RECT  4.350 0.615 4.510 0.715 ;
        RECT  3.385 0.275 4.440 0.365 ;
        RECT  4.260 0.455 4.350 0.715 ;
        RECT  3.730 0.455 4.260 0.545 ;
        RECT  4.070 0.635 4.170 0.745 ;
        RECT  4.070 1.120 4.125 1.525 ;
        RECT  3.980 0.635 4.070 1.525 ;
        RECT  3.350 1.055 3.980 1.165 ;
        RECT  3.620 0.455 3.730 0.935 ;
        RECT  3.275 0.275 3.385 0.535 ;
        RECT  3.265 1.255 3.375 1.525 ;
        RECT  3.260 0.625 3.350 1.165 ;
        RECT  3.050 0.445 3.275 0.535 ;
        RECT  3.150 1.255 3.265 1.345 ;
        RECT  3.160 0.625 3.260 0.725 ;
        RECT  3.060 0.820 3.150 1.345 ;
        RECT  1.915 1.435 3.140 1.525 ;
        RECT  2.870 0.265 3.130 0.355 ;
        RECT  3.050 0.820 3.060 0.910 ;
        RECT  2.960 0.445 3.050 0.910 ;
        RECT  2.760 0.265 2.870 0.365 ;
        RECT  0.665 0.275 2.760 0.365 ;
        RECT  2.560 1.215 2.675 1.325 ;
        RECT  2.560 0.455 2.625 0.800 ;
        RECT  2.515 0.455 2.560 1.325 ;
        RECT  2.470 0.700 2.515 1.325 ;
        RECT  1.945 0.700 2.470 0.800 ;
        RECT  1.230 0.495 2.395 0.585 ;
        RECT  1.235 1.205 2.380 1.315 ;
        RECT  1.855 0.700 1.945 1.095 ;
        RECT  1.705 1.405 1.915 1.525 ;
        RECT  1.340 1.000 1.855 1.095 ;
        RECT  0.635 1.435 1.705 1.525 ;
        RECT  0.900 0.725 1.290 0.835 ;
        RECT  0.785 0.470 0.900 1.345 ;
        RECT  0.400 0.990 0.785 1.100 ;
        RECT  0.475 0.275 0.665 0.405 ;
        RECT  0.525 1.270 0.635 1.525 ;
    END
END SDFXQD1

MACRO SDFXQD2
    CLASS CORE ;
    FOREIGN SDFXQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0583 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 0.890 ;
        RECT  0.430 0.670 0.450 0.890 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0650 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.000 2.950 1.290 ;
        RECT  2.780 1.000 2.850 1.090 ;
        RECT  2.650 0.910 2.780 1.090 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.865 0.565 6.950 1.150 ;
        RECT  6.850 0.275 6.865 1.460 ;
        RECT  6.760 0.275 6.850 0.665 ;
        RECT  6.760 1.050 6.850 1.460 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.890 2.350 1.090 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0322 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.890 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.850 4.350 1.290 ;
        RECT  4.160 0.850 4.250 1.020 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.125 -0.165 7.200 0.165 ;
        RECT  7.015 -0.165 7.125 0.485 ;
        RECT  4.790 -0.165 7.015 0.165 ;
        RECT  4.680 -0.165 4.790 0.420 ;
        RECT  0.185 -0.165 4.680 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.125 1.635 7.200 1.965 ;
        RECT  7.015 1.250 7.125 1.965 ;
        RECT  3.880 1.635 7.015 1.965 ;
        RECT  3.770 1.335 3.880 1.965 ;
        RECT  0.185 1.635 3.770 1.965 ;
        RECT  0.075 1.275 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.580 0.615 6.670 1.345 ;
        RECT  6.375 0.615 6.580 0.725 ;
        RECT  6.235 1.235 6.580 1.345 ;
        RECT  6.265 0.255 6.375 0.725 ;
        RECT  6.005 0.825 6.320 0.935 ;
        RECT  5.870 0.615 6.265 0.725 ;
        RECT  5.915 0.825 6.005 1.345 ;
        RECT  5.780 0.825 5.915 0.915 ;
        RECT  5.520 1.235 5.915 1.345 ;
        RECT  5.690 0.305 5.780 0.915 ;
        RECT  5.430 1.005 5.775 1.105 ;
        RECT  5.510 0.305 5.690 0.415 ;
        RECT  5.430 0.565 5.595 0.675 ;
        RECT  5.325 1.435 5.535 1.545 ;
        RECT  5.340 0.565 5.430 1.320 ;
        RECT  4.740 0.580 5.340 0.690 ;
        RECT  4.725 1.210 5.340 1.320 ;
        RECT  5.030 1.435 5.325 1.525 ;
        RECT  5.125 0.830 5.235 1.120 ;
        RECT  4.630 1.030 5.125 1.120 ;
        RECT  4.815 1.435 5.030 1.545 ;
        RECT  4.125 1.435 4.815 1.525 ;
        RECT  4.620 1.030 4.630 1.305 ;
        RECT  4.510 0.615 4.620 1.305 ;
        RECT  4.440 0.275 4.550 0.525 ;
        RECT  4.350 0.615 4.510 0.715 ;
        RECT  3.385 0.275 4.440 0.365 ;
        RECT  4.260 0.455 4.350 0.715 ;
        RECT  3.730 0.455 4.260 0.545 ;
        RECT  4.070 0.635 4.170 0.745 ;
        RECT  4.070 1.120 4.125 1.525 ;
        RECT  3.980 0.635 4.070 1.525 ;
        RECT  3.350 1.055 3.980 1.165 ;
        RECT  3.620 0.455 3.730 0.935 ;
        RECT  3.275 0.275 3.385 0.535 ;
        RECT  3.265 1.255 3.375 1.525 ;
        RECT  3.260 0.625 3.350 1.165 ;
        RECT  3.050 0.445 3.275 0.535 ;
        RECT  3.150 1.255 3.265 1.345 ;
        RECT  3.160 0.625 3.260 0.725 ;
        RECT  3.060 0.820 3.150 1.345 ;
        RECT  1.915 1.435 3.140 1.525 ;
        RECT  2.870 0.265 3.130 0.355 ;
        RECT  3.050 0.820 3.060 0.910 ;
        RECT  2.960 0.445 3.050 0.910 ;
        RECT  2.760 0.265 2.870 0.365 ;
        RECT  0.665 0.275 2.760 0.365 ;
        RECT  2.560 1.215 2.675 1.325 ;
        RECT  2.560 0.455 2.625 0.800 ;
        RECT  2.515 0.455 2.560 1.325 ;
        RECT  2.470 0.700 2.515 1.325 ;
        RECT  1.945 0.700 2.470 0.800 ;
        RECT  1.230 0.495 2.395 0.585 ;
        RECT  1.235 1.205 2.380 1.315 ;
        RECT  1.855 0.700 1.945 1.095 ;
        RECT  1.705 1.405 1.915 1.525 ;
        RECT  1.340 1.000 1.855 1.095 ;
        RECT  0.635 1.435 1.705 1.525 ;
        RECT  0.900 0.725 1.290 0.835 ;
        RECT  0.785 0.470 0.900 1.345 ;
        RECT  0.400 0.990 0.785 1.100 ;
        RECT  0.475 0.275 0.665 0.405 ;
        RECT  0.525 1.270 0.635 1.525 ;
    END
END SDFXQD2

MACRO SDFXQD4
    CLASS CORE ;
    FOREIGN SDFXQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0583 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 0.890 ;
        RECT  0.430 0.670 0.450 0.890 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0650 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.000 2.950 1.290 ;
        RECT  2.780 1.000 2.850 1.090 ;
        RECT  2.650 0.910 2.780 1.090 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 0.325 8.075 0.635 ;
        RECT  7.850 1.100 8.075 1.410 ;
        RECT  7.550 0.325 7.850 1.410 ;
        RECT  7.405 0.325 7.550 0.635 ;
        RECT  7.405 1.100 7.550 1.410 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.890 2.350 1.090 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0322 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.890 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0445 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.910 4.150 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.305 -0.165 8.400 0.165 ;
        RECT  8.195 -0.165 8.305 0.685 ;
        RECT  7.285 -0.165 8.195 0.165 ;
        RECT  7.175 -0.165 7.285 0.465 ;
        RECT  6.805 -0.165 7.175 0.165 ;
        RECT  6.635 -0.165 6.805 0.415 ;
        RECT  5.770 -0.165 6.635 0.165 ;
        RECT  5.600 -0.165 5.770 0.405 ;
        RECT  4.715 -0.165 5.600 0.165 ;
        RECT  4.605 -0.165 4.715 0.725 ;
        RECT  3.940 -0.165 4.605 0.165 ;
        RECT  3.770 -0.165 3.940 0.355 ;
        RECT  0.185 -0.165 3.770 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.305 1.635 8.400 1.965 ;
        RECT  8.195 1.050 8.305 1.965 ;
        RECT  5.880 1.635 8.195 1.965 ;
        RECT  5.790 1.135 5.880 1.965 ;
        RECT  5.625 1.135 5.790 1.245 ;
        RECT  0.185 1.635 5.790 1.965 ;
        RECT  0.075 1.275 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.950 0.325 8.075 0.635 ;
        RECT  7.950 1.100 8.075 1.410 ;
        RECT  7.405 0.325 7.450 0.635 ;
        RECT  7.405 1.100 7.450 1.410 ;
        RECT  7.105 0.585 7.195 1.495 ;
        RECT  7.040 0.585 7.105 0.675 ;
        RECT  6.895 1.385 7.105 1.495 ;
        RECT  6.920 0.275 7.040 0.675 ;
        RECT  6.715 0.780 7.005 0.890 ;
        RECT  6.645 0.585 6.920 0.675 ;
        RECT  6.610 0.780 6.715 1.495 ;
        RECT  6.535 0.505 6.645 0.675 ;
        RECT  6.420 0.780 6.610 0.890 ;
        RECT  6.060 1.385 6.610 1.495 ;
        RECT  6.240 1.120 6.490 1.230 ;
        RECT  6.330 0.305 6.420 0.890 ;
        RECT  5.965 0.305 6.330 0.415 ;
        RECT  6.190 0.735 6.240 1.230 ;
        RECT  6.150 0.560 6.190 1.230 ;
        RECT  6.080 0.560 6.150 0.845 ;
        RECT  4.975 0.735 6.080 0.845 ;
        RECT  5.970 0.955 6.060 1.495 ;
        RECT  5.480 0.955 5.970 1.045 ;
        RECT  5.875 0.305 5.965 0.605 ;
        RECT  5.235 0.495 5.875 0.605 ;
        RECT  5.480 1.345 5.700 1.515 ;
        RECT  5.370 0.955 5.480 1.165 ;
        RECT  5.370 1.255 5.480 1.515 ;
        RECT  5.185 1.055 5.370 1.165 ;
        RECT  4.705 1.255 5.370 1.345 ;
        RECT  5.065 1.435 5.240 1.545 ;
        RECT  5.125 0.335 5.235 0.605 ;
        RECT  4.975 1.055 5.095 1.165 ;
        RECT  4.375 1.435 5.065 1.525 ;
        RECT  4.865 0.490 4.975 1.165 ;
        RECT  4.580 1.175 4.705 1.345 ;
        RECT  4.480 1.175 4.580 1.285 ;
        RECT  4.165 0.305 4.480 0.415 ;
        RECT  4.390 0.515 4.480 1.285 ;
        RECT  4.345 0.515 4.390 0.725 ;
        RECT  3.760 1.180 4.390 1.285 ;
        RECT  4.245 1.385 4.375 1.525 ;
        RECT  3.560 1.385 4.245 1.495 ;
        RECT  3.560 0.625 4.225 0.735 ;
        RECT  4.075 0.305 4.165 0.535 ;
        RECT  3.445 0.445 4.075 0.535 ;
        RECT  3.670 0.915 3.760 1.285 ;
        RECT  3.470 0.625 3.560 1.495 ;
        RECT  3.175 0.625 3.470 0.735 ;
        RECT  3.420 1.075 3.470 1.245 ;
        RECT  3.315 0.275 3.445 0.535 ;
        RECT  3.310 1.355 3.365 1.525 ;
        RECT  3.085 0.445 3.315 0.535 ;
        RECT  3.210 0.825 3.310 1.525 ;
        RECT  3.085 0.825 3.210 0.915 ;
        RECT  2.865 0.265 3.130 0.355 ;
        RECT  3.005 1.365 3.115 1.545 ;
        RECT  2.995 0.445 3.085 0.915 ;
        RECT  1.915 1.435 3.005 1.525 ;
        RECT  2.760 0.265 2.865 0.365 ;
        RECT  0.665 0.275 2.760 0.365 ;
        RECT  2.560 1.215 2.675 1.325 ;
        RECT  2.560 0.455 2.625 0.800 ;
        RECT  2.515 0.455 2.560 1.325 ;
        RECT  2.470 0.700 2.515 1.325 ;
        RECT  1.945 0.700 2.470 0.800 ;
        RECT  1.230 0.495 2.395 0.585 ;
        RECT  1.235 1.205 2.380 1.315 ;
        RECT  1.855 0.700 1.945 1.095 ;
        RECT  1.705 1.405 1.915 1.525 ;
        RECT  1.340 1.000 1.855 1.095 ;
        RECT  0.635 1.435 1.705 1.525 ;
        RECT  0.900 0.725 1.290 0.835 ;
        RECT  0.785 0.470 0.900 1.345 ;
        RECT  0.400 0.990 0.785 1.100 ;
        RECT  0.475 0.275 0.665 0.405 ;
        RECT  0.525 1.270 0.635 1.525 ;
    END
END SDFXQD4

MACRO SEDFCND0
    CLASS CORE ;
    FOREIGN SEDFCND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0506 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.645 0.480 7.750 1.290 ;
        RECT  7.625 0.480 7.645 0.675 ;
        RECT  7.625 1.055 7.645 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.245 0.500 7.355 1.170 ;
        RECT  7.110 0.500 7.245 0.690 ;
        RECT  7.070 1.060 7.245 1.170 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0662 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0219 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.510 3.355 0.895 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0575 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.645 0.480 6.755 1.000 ;
        RECT  6.450 0.890 6.645 1.000 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.180 -0.165 7.800 0.165 ;
        RECT  6.010 -0.165 6.180 0.355 ;
        RECT  4.940 -0.165 6.010 0.165 ;
        RECT  4.830 -0.165 4.940 0.405 ;
        RECT  0.185 -0.165 4.830 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.470 1.635 7.800 1.965 ;
        RECT  7.300 1.505 7.470 1.965 ;
        RECT  7.020 1.635 7.300 1.965 ;
        RECT  6.850 1.505 7.020 1.965 ;
        RECT  5.220 1.635 6.850 1.965 ;
        RECT  5.050 1.445 5.220 1.965 ;
        RECT  0.185 1.635 5.050 1.965 ;
        RECT  0.075 1.300 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.535 0.775 7.555 0.945 ;
        RECT  7.445 0.775 7.535 1.415 ;
        RECT  6.160 1.325 7.445 1.415 ;
        RECT  6.970 0.780 7.135 0.890 ;
        RECT  6.960 0.460 6.970 0.890 ;
        RECT  6.850 0.460 6.960 1.235 ;
        RECT  6.535 0.275 6.935 0.365 ;
        RECT  6.300 1.130 6.850 1.235 ;
        RECT  6.445 0.275 6.535 0.535 ;
        RECT  5.850 0.445 6.445 0.535 ;
        RECT  6.190 0.860 6.300 1.235 ;
        RECT  6.075 0.625 6.255 0.735 ;
        RECT  6.075 1.325 6.160 1.515 ;
        RECT  5.985 0.625 6.075 1.515 ;
        RECT  5.965 0.625 5.985 0.785 ;
        RECT  5.410 1.425 5.985 1.515 ;
        RECT  5.755 0.685 5.965 0.785 ;
        RECT  5.765 0.875 5.875 1.335 ;
        RECT  5.740 0.445 5.850 0.595 ;
        RECT  5.645 0.875 5.765 0.975 ;
        RECT  5.645 0.505 5.740 0.595 ;
        RECT  5.530 0.505 5.645 0.975 ;
        RECT  5.505 1.065 5.615 1.315 ;
        RECT  5.120 0.305 5.550 0.415 ;
        RECT  5.430 1.065 5.505 1.155 ;
        RECT  5.340 0.505 5.430 1.155 ;
        RECT  5.310 1.265 5.410 1.515 ;
        RECT  5.210 0.505 5.340 0.615 ;
        RECT  4.590 0.905 5.340 0.995 ;
        RECT  4.960 1.265 5.310 1.355 ;
        RECT  4.300 0.705 5.240 0.815 ;
        RECT  4.780 1.085 5.180 1.175 ;
        RECT  5.030 0.305 5.120 0.585 ;
        RECT  4.690 0.495 5.030 0.585 ;
        RECT  4.870 1.265 4.960 1.525 ;
        RECT  4.055 1.435 4.870 1.525 ;
        RECT  4.680 1.085 4.780 1.255 ;
        RECT  4.600 0.305 4.690 0.585 ;
        RECT  4.480 1.145 4.680 1.255 ;
        RECT  4.180 0.305 4.600 0.415 ;
        RECT  4.420 0.905 4.590 1.015 ;
        RECT  4.185 0.525 4.300 1.325 ;
        RECT  4.060 0.525 4.185 0.635 ;
        RECT  3.940 0.915 4.080 1.025 ;
        RECT  3.965 1.255 4.055 1.525 ;
        RECT  2.575 1.255 3.965 1.345 ;
        RECT  3.750 0.275 3.960 0.385 ;
        RECT  3.840 0.520 3.940 1.165 ;
        RECT  3.700 1.435 3.875 1.545 ;
        RECT  3.525 0.520 3.840 0.630 ;
        RECT  3.625 1.055 3.840 1.165 ;
        RECT  0.710 0.275 3.750 0.365 ;
        RECT  3.535 0.750 3.740 0.860 ;
        RECT  1.955 1.435 3.700 1.525 ;
        RECT  3.445 0.750 3.535 1.165 ;
        RECT  3.150 1.055 3.445 1.165 ;
        RECT  3.040 0.490 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.675 2.755 1.165 ;
        RECT  2.665 0.495 2.670 1.165 ;
        RECT  2.560 0.495 2.665 0.765 ;
        RECT  2.485 0.890 2.575 1.345 ;
        RECT  2.055 0.675 2.560 0.765 ;
        RECT  2.170 0.890 2.485 1.000 ;
        RECT  1.215 0.475 2.435 0.585 ;
        RECT  2.285 1.130 2.395 1.305 ;
        RECT  1.455 1.215 2.285 1.305 ;
        RECT  1.945 0.675 2.055 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.945 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.330 1.005 1.520 1.125 ;
        RECT  1.245 1.215 1.455 1.345 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.905 0.510 0.910 0.835 ;
        RECT  0.795 0.510 0.905 1.345 ;
        RECT  0.720 0.510 0.795 0.620 ;
        RECT  0.410 0.990 0.795 1.100 ;
        RECT  0.500 0.255 0.710 0.365 ;
        RECT  0.535 1.300 0.645 1.525 ;
    END
END SEDFCND0

MACRO SEDFCND1
    CLASS CORE ;
    FOREIGN SEDFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0569 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.645 0.275 7.750 1.490 ;
        RECT  7.615 0.275 7.645 0.675 ;
        RECT  7.625 1.050 7.645 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.245 0.565 7.355 1.170 ;
        RECT  7.220 0.565 7.245 0.665 ;
        RECT  7.070 1.060 7.245 1.170 ;
        RECT  7.110 0.275 7.220 0.665 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0725 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.510 3.355 0.895 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0575 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.645 0.480 6.755 1.000 ;
        RECT  6.450 0.890 6.645 1.000 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.180 -0.165 7.800 0.165 ;
        RECT  6.010 -0.165 6.180 0.355 ;
        RECT  4.940 -0.165 6.010 0.165 ;
        RECT  4.830 -0.165 4.940 0.405 ;
        RECT  0.185 -0.165 4.830 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.020 1.635 7.800 1.965 ;
        RECT  6.850 1.505 7.020 1.965 ;
        RECT  5.220 1.635 6.850 1.965 ;
        RECT  5.050 1.445 5.220 1.965 ;
        RECT  0.185 1.635 5.050 1.965 ;
        RECT  0.075 1.300 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.535 0.775 7.555 0.945 ;
        RECT  7.445 0.775 7.535 1.415 ;
        RECT  6.160 1.325 7.445 1.415 ;
        RECT  6.970 0.780 7.135 0.890 ;
        RECT  6.960 0.460 6.970 0.890 ;
        RECT  6.850 0.460 6.960 1.235 ;
        RECT  6.535 0.275 6.935 0.365 ;
        RECT  6.300 1.130 6.850 1.235 ;
        RECT  6.445 0.275 6.535 0.535 ;
        RECT  5.850 0.445 6.445 0.535 ;
        RECT  6.190 0.860 6.300 1.235 ;
        RECT  6.075 0.625 6.255 0.735 ;
        RECT  6.075 1.325 6.160 1.515 ;
        RECT  5.985 0.625 6.075 1.515 ;
        RECT  5.965 0.625 5.985 0.785 ;
        RECT  5.410 1.425 5.985 1.515 ;
        RECT  5.755 0.685 5.965 0.785 ;
        RECT  5.765 0.875 5.875 1.335 ;
        RECT  5.740 0.445 5.850 0.595 ;
        RECT  5.645 0.875 5.765 0.975 ;
        RECT  5.645 0.505 5.740 0.595 ;
        RECT  5.530 0.505 5.645 0.975 ;
        RECT  5.505 1.065 5.615 1.315 ;
        RECT  5.120 0.305 5.550 0.415 ;
        RECT  5.430 1.065 5.505 1.155 ;
        RECT  5.340 0.505 5.430 1.155 ;
        RECT  5.310 1.265 5.410 1.515 ;
        RECT  5.210 0.505 5.340 0.615 ;
        RECT  4.590 0.905 5.340 0.995 ;
        RECT  4.960 1.265 5.310 1.355 ;
        RECT  4.300 0.705 5.240 0.815 ;
        RECT  4.780 1.085 5.180 1.175 ;
        RECT  5.030 0.305 5.120 0.585 ;
        RECT  4.690 0.495 5.030 0.585 ;
        RECT  4.870 1.265 4.960 1.525 ;
        RECT  4.055 1.435 4.870 1.525 ;
        RECT  4.680 1.085 4.780 1.255 ;
        RECT  4.600 0.305 4.690 0.585 ;
        RECT  4.480 1.145 4.680 1.255 ;
        RECT  4.180 0.305 4.600 0.415 ;
        RECT  4.420 0.905 4.590 1.015 ;
        RECT  4.185 0.525 4.300 1.325 ;
        RECT  4.060 0.525 4.185 0.635 ;
        RECT  3.940 0.915 4.080 1.025 ;
        RECT  3.965 1.255 4.055 1.525 ;
        RECT  2.575 1.255 3.965 1.345 ;
        RECT  3.750 0.275 3.960 0.385 ;
        RECT  3.840 0.520 3.940 1.165 ;
        RECT  3.700 1.435 3.875 1.545 ;
        RECT  3.525 0.520 3.840 0.630 ;
        RECT  3.625 1.055 3.840 1.165 ;
        RECT  0.710 0.275 3.750 0.365 ;
        RECT  3.535 0.750 3.740 0.860 ;
        RECT  1.955 1.435 3.700 1.525 ;
        RECT  3.445 0.750 3.535 1.165 ;
        RECT  3.150 1.055 3.445 1.165 ;
        RECT  3.040 0.455 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.675 2.755 1.165 ;
        RECT  2.665 0.475 2.670 1.165 ;
        RECT  2.560 0.475 2.665 0.765 ;
        RECT  2.485 0.890 2.575 1.345 ;
        RECT  2.055 0.675 2.560 0.765 ;
        RECT  2.170 0.890 2.485 1.000 ;
        RECT  1.215 0.475 2.435 0.585 ;
        RECT  2.285 1.130 2.395 1.305 ;
        RECT  1.455 1.215 2.285 1.305 ;
        RECT  1.945 0.675 2.055 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.945 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.330 1.005 1.520 1.125 ;
        RECT  1.245 1.215 1.455 1.345 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.795 0.510 0.910 1.345 ;
        RECT  0.720 0.510 0.795 0.620 ;
        RECT  0.410 0.990 0.795 1.100 ;
        RECT  0.500 0.255 0.710 0.365 ;
        RECT  0.535 1.300 0.645 1.525 ;
    END
END SEDFCND1

MACRO SEDFCND2
    CLASS CORE ;
    FOREIGN SEDFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0569 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 0.285 7.950 1.490 ;
        RECT  7.765 0.285 7.850 0.665 ;
        RECT  7.765 1.075 7.850 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.240 0.285 7.375 1.240 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0725 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.510 3.355 0.895 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0575 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.510 6.550 1.030 ;
        RECT  6.440 0.820 6.450 1.030 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.180 -0.165 8.200 0.165 ;
        RECT  6.010 -0.165 6.180 0.355 ;
        RECT  4.940 -0.165 6.010 0.165 ;
        RECT  4.830 -0.165 4.940 0.405 ;
        RECT  0.185 -0.165 4.830 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.060 1.635 8.200 1.965 ;
        RECT  6.890 1.515 7.060 1.965 ;
        RECT  5.220 1.635 6.890 1.965 ;
        RECT  5.050 1.445 5.220 1.965 ;
        RECT  0.185 1.635 5.050 1.965 ;
        RECT  0.075 1.300 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.620 0.780 7.760 0.890 ;
        RECT  7.530 0.780 7.620 1.425 ;
        RECT  6.075 1.330 7.530 1.425 ;
        RECT  7.020 0.510 7.130 1.240 ;
        RECT  6.735 0.510 7.020 0.620 ;
        RECT  6.300 1.130 7.020 1.240 ;
        RECT  6.360 0.275 6.875 0.375 ;
        RECT  6.270 0.275 6.360 0.535 ;
        RECT  6.190 0.860 6.300 1.240 ;
        RECT  5.850 0.445 6.270 0.535 ;
        RECT  6.075 0.625 6.255 0.735 ;
        RECT  5.985 0.625 6.075 1.515 ;
        RECT  5.965 0.625 5.985 0.785 ;
        RECT  5.410 1.425 5.985 1.515 ;
        RECT  5.755 0.685 5.965 0.785 ;
        RECT  5.765 0.875 5.875 1.335 ;
        RECT  5.740 0.445 5.850 0.595 ;
        RECT  5.645 0.875 5.765 0.975 ;
        RECT  5.645 0.505 5.740 0.595 ;
        RECT  5.530 0.505 5.645 0.975 ;
        RECT  5.505 1.065 5.615 1.315 ;
        RECT  5.120 0.305 5.550 0.415 ;
        RECT  5.430 1.065 5.505 1.155 ;
        RECT  5.340 0.505 5.430 1.155 ;
        RECT  5.310 1.265 5.410 1.515 ;
        RECT  5.210 0.505 5.340 0.615 ;
        RECT  4.590 0.905 5.340 0.995 ;
        RECT  4.960 1.265 5.310 1.355 ;
        RECT  4.300 0.705 5.240 0.815 ;
        RECT  4.780 1.085 5.180 1.175 ;
        RECT  5.030 0.305 5.120 0.585 ;
        RECT  4.690 0.495 5.030 0.585 ;
        RECT  4.870 1.265 4.960 1.525 ;
        RECT  4.055 1.435 4.870 1.525 ;
        RECT  4.680 1.085 4.780 1.255 ;
        RECT  4.600 0.305 4.690 0.585 ;
        RECT  4.480 1.145 4.680 1.255 ;
        RECT  4.180 0.305 4.600 0.415 ;
        RECT  4.420 0.905 4.590 1.015 ;
        RECT  4.185 0.525 4.300 1.325 ;
        RECT  4.060 0.525 4.185 0.635 ;
        RECT  3.940 0.915 4.080 1.025 ;
        RECT  3.965 1.255 4.055 1.525 ;
        RECT  2.575 1.255 3.965 1.345 ;
        RECT  3.750 0.275 3.960 0.385 ;
        RECT  3.840 0.520 3.940 1.165 ;
        RECT  3.700 1.435 3.875 1.545 ;
        RECT  3.525 0.520 3.840 0.630 ;
        RECT  3.625 1.055 3.840 1.165 ;
        RECT  0.710 0.275 3.750 0.365 ;
        RECT  3.535 0.750 3.740 0.860 ;
        RECT  1.955 1.435 3.700 1.525 ;
        RECT  3.445 0.750 3.535 1.165 ;
        RECT  3.150 1.055 3.445 1.165 ;
        RECT  3.040 0.455 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.675 2.755 1.165 ;
        RECT  2.665 0.475 2.670 1.165 ;
        RECT  2.560 0.475 2.665 0.765 ;
        RECT  2.485 0.890 2.575 1.345 ;
        RECT  2.055 0.675 2.560 0.765 ;
        RECT  2.170 0.890 2.485 1.000 ;
        RECT  1.215 0.475 2.435 0.585 ;
        RECT  2.285 1.130 2.395 1.305 ;
        RECT  1.455 1.215 2.285 1.305 ;
        RECT  1.945 0.675 2.055 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.945 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.330 1.005 1.520 1.125 ;
        RECT  1.245 1.215 1.455 1.345 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.795 0.510 0.910 1.345 ;
        RECT  0.720 0.510 0.795 0.620 ;
        RECT  0.410 0.990 0.795 1.100 ;
        RECT  0.500 0.255 0.710 0.365 ;
        RECT  0.535 1.300 0.645 1.525 ;
    END
END SEDFCND2

MACRO SEDFCND4
    CLASS CORE ;
    FOREIGN SEDFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0569 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.250 0.325 9.495 0.635 ;
        RECT  9.250 1.100 9.495 1.410 ;
        RECT  8.950 0.325 9.250 1.410 ;
        RECT  8.825 0.325 8.950 0.635 ;
        RECT  8.825 1.100 8.950 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.250 0.325 8.475 0.635 ;
        RECT  8.250 1.110 8.475 1.290 ;
        RECT  7.950 0.325 8.250 1.290 ;
        RECT  7.805 0.325 7.950 0.635 ;
        RECT  7.805 1.110 7.950 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0724 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.465 3.355 0.905 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1088 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.710 7.150 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.725 -0.165 9.800 0.165 ;
        RECT  9.615 -0.165 9.725 0.675 ;
        RECT  8.705 -0.165 9.615 0.165 ;
        RECT  8.595 -0.165 8.705 0.675 ;
        RECT  7.715 -0.165 8.595 0.165 ;
        RECT  7.520 -0.165 7.715 0.420 ;
        RECT  6.630 -0.165 7.520 0.165 ;
        RECT  6.440 -0.165 6.630 0.400 ;
        RECT  4.995 -0.165 6.440 0.165 ;
        RECT  4.885 -0.165 4.995 0.405 ;
        RECT  0.185 -0.165 4.885 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.725 1.635 9.800 1.965 ;
        RECT  9.615 1.050 9.725 1.965 ;
        RECT  5.275 1.635 9.615 1.965 ;
        RECT  5.105 1.445 5.275 1.965 ;
        RECT  0.185 1.635 5.105 1.965 ;
        RECT  0.075 1.285 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.350 0.325 9.495 0.635 ;
        RECT  9.350 1.100 9.495 1.410 ;
        RECT  8.825 0.325 8.850 0.635 ;
        RECT  8.825 1.100 8.850 1.410 ;
        RECT  8.350 0.325 8.475 0.635 ;
        RECT  8.350 1.110 8.475 1.290 ;
        RECT  7.805 0.325 7.850 0.635 ;
        RECT  7.805 1.110 7.850 1.290 ;
        RECT  8.710 0.790 8.825 0.900 ;
        RECT  8.620 0.790 8.710 1.515 ;
        RECT  6.245 1.425 8.620 1.515 ;
        RECT  7.670 0.785 7.830 0.895 ;
        RECT  7.580 0.510 7.670 1.285 ;
        RECT  6.560 0.510 7.580 0.600 ;
        RECT  6.715 1.175 7.580 1.285 ;
        RECT  7.380 0.730 7.490 1.070 ;
        RECT  6.760 0.980 7.380 1.070 ;
        RECT  6.660 0.710 6.760 1.070 ;
        RECT  6.565 0.980 6.660 1.070 ;
        RECT  6.440 0.980 6.565 1.305 ;
        RECT  6.450 0.510 6.560 0.865 ;
        RECT  6.260 0.755 6.450 0.865 ;
        RECT  5.930 1.215 6.440 1.305 ;
        RECT  6.165 0.505 6.335 0.615 ;
        RECT  6.165 1.015 6.265 1.125 ;
        RECT  6.075 1.395 6.245 1.515 ;
        RECT  5.175 0.305 6.195 0.415 ;
        RECT  6.075 0.505 6.165 1.125 ;
        RECT  5.820 0.505 6.075 0.615 ;
        RECT  5.465 1.425 6.075 1.515 ;
        RECT  5.820 0.865 5.930 1.305 ;
        RECT  5.700 0.865 5.820 0.975 ;
        RECT  5.585 0.515 5.700 0.975 ;
        RECT  5.560 1.065 5.670 1.315 ;
        RECT  5.485 1.065 5.560 1.155 ;
        RECT  5.395 0.505 5.485 1.155 ;
        RECT  5.365 1.265 5.465 1.515 ;
        RECT  5.265 0.505 5.395 0.615 ;
        RECT  4.635 0.905 5.395 0.995 ;
        RECT  5.015 1.265 5.365 1.355 ;
        RECT  4.455 0.705 5.295 0.815 ;
        RECT  4.835 1.085 5.235 1.175 ;
        RECT  5.085 0.305 5.175 0.585 ;
        RECT  4.745 0.495 5.085 0.585 ;
        RECT  4.925 1.265 5.015 1.525 ;
        RECT  4.345 1.435 4.925 1.525 ;
        RECT  4.725 1.085 4.835 1.310 ;
        RECT  4.655 0.305 4.745 0.585 ;
        RECT  4.535 1.200 4.725 1.310 ;
        RECT  4.175 0.305 4.655 0.415 ;
        RECT  4.545 0.905 4.635 1.090 ;
        RECT  4.365 0.525 4.455 1.125 ;
        RECT  4.095 0.525 4.365 0.635 ;
        RECT  4.220 1.015 4.365 1.125 ;
        RECT  4.235 1.255 4.345 1.525 ;
        RECT  4.165 0.740 4.275 0.910 ;
        RECT  2.575 1.255 4.235 1.345 ;
        RECT  3.965 0.800 4.165 0.910 ;
        RECT  3.900 1.435 4.095 1.545 ;
        RECT  3.560 0.275 3.965 0.385 ;
        RECT  3.855 0.520 3.965 1.165 ;
        RECT  1.955 1.435 3.900 1.525 ;
        RECT  3.560 0.520 3.855 0.630 ;
        RECT  3.625 1.045 3.855 1.165 ;
        RECT  3.535 0.780 3.655 0.890 ;
        RECT  0.690 0.275 3.560 0.365 ;
        RECT  3.445 0.780 3.535 1.165 ;
        RECT  3.150 1.045 3.445 1.165 ;
        RECT  3.040 0.455 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.710 2.755 1.165 ;
        RECT  2.665 0.490 2.670 1.165 ;
        RECT  2.560 0.490 2.665 0.800 ;
        RECT  2.485 0.900 2.575 1.345 ;
        RECT  2.065 0.710 2.560 0.800 ;
        RECT  2.170 0.900 2.485 1.010 ;
        RECT  1.210 0.475 2.435 0.585 ;
        RECT  2.280 1.130 2.395 1.305 ;
        RECT  1.600 1.215 2.280 1.305 ;
        RECT  1.935 0.675 2.065 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.935 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.245 1.215 1.600 1.345 ;
        RECT  1.330 1.015 1.520 1.125 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.795 0.520 0.910 1.345 ;
        RECT  0.720 0.520 0.795 0.610 ;
        RECT  0.400 1.000 0.795 1.090 ;
        RECT  0.475 0.265 0.690 0.365 ;
        RECT  0.535 1.300 0.645 1.525 ;
    END
END SEDFCND4

MACRO SEDFCNQD0
    CLASS CORE ;
    FOREIGN SEDFCNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0506 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.265 0.590 7.355 1.170 ;
        RECT  7.245 0.280 7.265 1.480 ;
        RECT  7.155 0.280 7.245 0.690 ;
        RECT  7.155 1.060 7.245 1.480 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0559 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0219 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.510 3.355 0.895 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0575 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.645 0.480 6.755 1.000 ;
        RECT  6.450 0.890 6.645 1.000 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.525 -0.165 7.600 0.165 ;
        RECT  7.415 -0.165 7.525 0.480 ;
        RECT  6.180 -0.165 7.415 0.165 ;
        RECT  6.010 -0.165 6.180 0.355 ;
        RECT  4.940 -0.165 6.010 0.165 ;
        RECT  4.830 -0.165 4.940 0.405 ;
        RECT  0.185 -0.165 4.830 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.525 1.635 7.600 1.965 ;
        RECT  7.415 1.275 7.525 1.965 ;
        RECT  6.990 1.635 7.415 1.965 ;
        RECT  6.880 1.345 6.990 1.965 ;
        RECT  6.435 1.635 6.880 1.965 ;
        RECT  6.325 1.345 6.435 1.965 ;
        RECT  5.220 1.635 6.325 1.965 ;
        RECT  5.050 1.445 5.220 1.965 ;
        RECT  0.185 1.635 5.050 1.965 ;
        RECT  0.075 1.300 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.960 0.815 7.135 0.925 ;
        RECT  6.850 0.460 6.960 1.235 ;
        RECT  6.535 0.275 6.935 0.365 ;
        RECT  6.705 1.130 6.850 1.235 ;
        RECT  6.595 1.130 6.705 1.500 ;
        RECT  6.300 1.130 6.595 1.235 ;
        RECT  6.445 0.275 6.535 0.535 ;
        RECT  5.850 0.445 6.445 0.535 ;
        RECT  6.190 0.860 6.300 1.235 ;
        RECT  6.075 0.625 6.255 0.735 ;
        RECT  6.075 1.325 6.190 1.435 ;
        RECT  5.985 0.625 6.075 1.515 ;
        RECT  5.965 0.625 5.985 0.785 ;
        RECT  5.410 1.425 5.985 1.515 ;
        RECT  5.755 0.685 5.965 0.785 ;
        RECT  5.765 0.875 5.875 1.335 ;
        RECT  5.740 0.445 5.850 0.595 ;
        RECT  5.645 0.875 5.765 0.975 ;
        RECT  5.645 0.505 5.740 0.595 ;
        RECT  5.530 0.505 5.645 0.975 ;
        RECT  5.505 1.065 5.615 1.315 ;
        RECT  5.120 0.305 5.550 0.415 ;
        RECT  5.430 1.065 5.505 1.155 ;
        RECT  5.340 0.505 5.430 1.155 ;
        RECT  5.310 1.265 5.410 1.515 ;
        RECT  5.210 0.505 5.340 0.615 ;
        RECT  4.590 0.905 5.340 0.995 ;
        RECT  4.960 1.265 5.310 1.355 ;
        RECT  4.300 0.705 5.240 0.815 ;
        RECT  4.780 1.085 5.180 1.175 ;
        RECT  5.030 0.305 5.120 0.585 ;
        RECT  4.690 0.495 5.030 0.585 ;
        RECT  4.870 1.265 4.960 1.525 ;
        RECT  4.055 1.435 4.870 1.525 ;
        RECT  4.680 1.085 4.780 1.255 ;
        RECT  4.600 0.305 4.690 0.585 ;
        RECT  4.480 1.145 4.680 1.255 ;
        RECT  4.180 0.305 4.600 0.415 ;
        RECT  4.420 0.905 4.590 1.015 ;
        RECT  4.185 0.525 4.300 1.325 ;
        RECT  4.060 0.525 4.185 0.635 ;
        RECT  3.940 0.915 4.080 1.025 ;
        RECT  3.965 1.255 4.055 1.525 ;
        RECT  2.575 1.255 3.965 1.345 ;
        RECT  3.750 0.275 3.960 0.385 ;
        RECT  3.840 0.520 3.940 1.165 ;
        RECT  3.700 1.435 3.875 1.545 ;
        RECT  3.525 0.520 3.840 0.630 ;
        RECT  3.625 1.055 3.840 1.165 ;
        RECT  0.710 0.275 3.750 0.365 ;
        RECT  3.535 0.750 3.740 0.860 ;
        RECT  1.955 1.435 3.700 1.525 ;
        RECT  3.445 0.750 3.535 1.165 ;
        RECT  3.150 1.055 3.445 1.165 ;
        RECT  3.040 0.490 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.675 2.755 1.165 ;
        RECT  2.665 0.495 2.670 1.165 ;
        RECT  2.560 0.495 2.665 0.765 ;
        RECT  2.485 0.890 2.575 1.345 ;
        RECT  2.055 0.675 2.560 0.765 ;
        RECT  2.170 0.890 2.485 1.000 ;
        RECT  1.215 0.475 2.435 0.585 ;
        RECT  2.285 1.130 2.395 1.305 ;
        RECT  1.455 1.215 2.285 1.305 ;
        RECT  1.945 0.675 2.055 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.945 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.330 1.005 1.520 1.125 ;
        RECT  1.245 1.215 1.455 1.345 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.905 0.510 0.910 0.835 ;
        RECT  0.795 0.510 0.905 1.345 ;
        RECT  0.720 0.510 0.795 0.620 ;
        RECT  0.410 0.990 0.795 1.100 ;
        RECT  0.500 0.255 0.710 0.365 ;
        RECT  0.535 1.300 0.645 1.525 ;
    END
END SEDFCNQD0

MACRO SEDFCNQD1
    CLASS CORE ;
    FOREIGN SEDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0569 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1560 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.265 0.590 7.355 1.170 ;
        RECT  7.245 0.280 7.265 1.480 ;
        RECT  7.155 0.280 7.245 0.690 ;
        RECT  7.155 1.060 7.245 1.480 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0725 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.510 3.355 0.895 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0575 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.645 0.480 6.755 1.000 ;
        RECT  6.450 0.890 6.645 1.000 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.525 -0.165 7.600 0.165 ;
        RECT  7.415 -0.165 7.525 0.480 ;
        RECT  6.180 -0.165 7.415 0.165 ;
        RECT  6.010 -0.165 6.180 0.355 ;
        RECT  4.940 -0.165 6.010 0.165 ;
        RECT  4.830 -0.165 4.940 0.405 ;
        RECT  0.185 -0.165 4.830 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.525 1.635 7.600 1.965 ;
        RECT  7.415 1.275 7.525 1.965 ;
        RECT  6.990 1.635 7.415 1.965 ;
        RECT  6.880 1.345 6.990 1.965 ;
        RECT  6.435 1.635 6.880 1.965 ;
        RECT  6.325 1.345 6.435 1.965 ;
        RECT  5.220 1.635 6.325 1.965 ;
        RECT  5.050 1.445 5.220 1.965 ;
        RECT  0.185 1.635 5.050 1.965 ;
        RECT  0.075 1.300 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.960 0.780 7.135 0.890 ;
        RECT  6.850 0.460 6.960 1.225 ;
        RECT  6.535 0.275 6.935 0.365 ;
        RECT  6.705 1.130 6.850 1.225 ;
        RECT  6.595 1.130 6.705 1.500 ;
        RECT  6.300 1.130 6.595 1.225 ;
        RECT  6.445 0.275 6.535 0.535 ;
        RECT  5.850 0.445 6.445 0.535 ;
        RECT  6.190 0.860 6.300 1.225 ;
        RECT  6.075 0.625 6.255 0.735 ;
        RECT  6.075 1.315 6.190 1.425 ;
        RECT  5.985 0.625 6.075 1.515 ;
        RECT  5.965 0.625 5.985 0.785 ;
        RECT  5.410 1.425 5.985 1.515 ;
        RECT  5.755 0.685 5.965 0.785 ;
        RECT  5.765 0.875 5.875 1.335 ;
        RECT  5.740 0.445 5.850 0.595 ;
        RECT  5.645 0.875 5.765 0.975 ;
        RECT  5.645 0.505 5.740 0.595 ;
        RECT  5.530 0.505 5.645 0.975 ;
        RECT  5.505 1.065 5.615 1.315 ;
        RECT  5.120 0.305 5.550 0.415 ;
        RECT  5.430 1.065 5.505 1.155 ;
        RECT  5.340 0.505 5.430 1.155 ;
        RECT  5.310 1.265 5.410 1.515 ;
        RECT  5.210 0.505 5.340 0.615 ;
        RECT  4.590 0.905 5.340 0.995 ;
        RECT  4.960 1.265 5.310 1.355 ;
        RECT  4.300 0.705 5.240 0.815 ;
        RECT  4.780 1.085 5.180 1.175 ;
        RECT  5.030 0.305 5.120 0.585 ;
        RECT  4.690 0.495 5.030 0.585 ;
        RECT  4.870 1.265 4.960 1.525 ;
        RECT  4.055 1.435 4.870 1.525 ;
        RECT  4.680 1.085 4.780 1.255 ;
        RECT  4.600 0.305 4.690 0.585 ;
        RECT  4.480 1.145 4.680 1.255 ;
        RECT  4.180 0.305 4.600 0.415 ;
        RECT  4.420 0.905 4.590 1.015 ;
        RECT  4.185 0.525 4.300 1.325 ;
        RECT  4.060 0.525 4.185 0.635 ;
        RECT  3.940 0.915 4.080 1.025 ;
        RECT  3.965 1.255 4.055 1.525 ;
        RECT  2.575 1.255 3.965 1.345 ;
        RECT  3.750 0.275 3.960 0.385 ;
        RECT  3.840 0.520 3.940 1.165 ;
        RECT  3.700 1.435 3.875 1.545 ;
        RECT  3.525 0.520 3.840 0.630 ;
        RECT  3.625 1.055 3.840 1.165 ;
        RECT  0.710 0.275 3.750 0.365 ;
        RECT  3.535 0.750 3.740 0.860 ;
        RECT  1.955 1.435 3.700 1.525 ;
        RECT  3.445 0.750 3.535 1.165 ;
        RECT  3.150 1.055 3.445 1.165 ;
        RECT  3.040 0.455 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.675 2.755 1.165 ;
        RECT  2.665 0.475 2.670 1.165 ;
        RECT  2.560 0.475 2.665 0.765 ;
        RECT  2.485 0.890 2.575 1.345 ;
        RECT  2.055 0.675 2.560 0.765 ;
        RECT  2.170 0.890 2.485 1.000 ;
        RECT  1.215 0.475 2.435 0.585 ;
        RECT  2.285 1.130 2.395 1.305 ;
        RECT  1.455 1.215 2.285 1.305 ;
        RECT  1.945 0.675 2.055 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.945 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.330 1.005 1.520 1.125 ;
        RECT  1.245 1.215 1.455 1.345 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.795 0.510 0.910 1.345 ;
        RECT  0.720 0.510 0.795 0.620 ;
        RECT  0.410 0.990 0.795 1.100 ;
        RECT  0.500 0.255 0.710 0.365 ;
        RECT  0.535 1.300 0.645 1.525 ;
    END
END SEDFCNQD1

MACRO SEDFCNQD2
    CLASS CORE ;
    FOREIGN SEDFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0593 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.475 0.590 7.555 1.170 ;
        RECT  7.445 0.280 7.475 1.480 ;
        RECT  7.345 0.280 7.445 0.690 ;
        RECT  7.350 1.060 7.445 1.480 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0725 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.510 3.355 0.895 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0575 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.630 0.480 6.755 1.000 ;
        RECT  6.435 0.890 6.630 1.000 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.735 -0.165 7.800 0.165 ;
        RECT  7.605 -0.165 7.735 0.480 ;
        RECT  7.215 -0.165 7.605 0.165 ;
        RECT  7.090 -0.165 7.215 0.690 ;
        RECT  6.180 -0.165 7.090 0.165 ;
        RECT  6.010 -0.165 6.180 0.355 ;
        RECT  4.940 -0.165 6.010 0.165 ;
        RECT  4.830 -0.165 4.940 0.405 ;
        RECT  0.185 -0.165 4.830 0.165 ;
        RECT  0.075 -0.165 0.185 0.495 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.735 1.635 7.800 1.965 ;
        RECT  7.605 1.275 7.735 1.965 ;
        RECT  7.215 1.635 7.605 1.965 ;
        RECT  7.085 1.020 7.215 1.965 ;
        RECT  6.815 1.375 7.085 1.485 ;
        RECT  6.470 1.635 7.085 1.965 ;
        RECT  6.285 1.370 6.470 1.965 ;
        RECT  5.220 1.635 6.285 1.965 ;
        RECT  5.050 1.445 5.220 1.965 ;
        RECT  0.185 1.635 5.050 1.965 ;
        RECT  0.075 1.220 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.960 0.815 7.335 0.925 ;
        RECT  6.845 0.475 6.960 1.280 ;
        RECT  6.465 0.275 6.920 0.365 ;
        RECT  6.300 1.160 6.845 1.280 ;
        RECT  6.375 0.275 6.465 0.535 ;
        RECT  5.850 0.445 6.375 0.535 ;
        RECT  6.190 0.860 6.300 1.280 ;
        RECT  6.075 0.625 6.255 0.735 ;
        RECT  6.075 1.370 6.195 1.515 ;
        RECT  5.985 0.625 6.075 1.515 ;
        RECT  5.965 0.625 5.985 0.775 ;
        RECT  5.410 1.425 5.985 1.515 ;
        RECT  5.755 0.685 5.965 0.775 ;
        RECT  5.765 0.865 5.875 1.335 ;
        RECT  5.740 0.445 5.850 0.595 ;
        RECT  5.645 0.865 5.765 0.975 ;
        RECT  5.645 0.505 5.740 0.595 ;
        RECT  5.530 0.505 5.645 0.975 ;
        RECT  5.505 1.065 5.615 1.315 ;
        RECT  5.120 0.305 5.550 0.415 ;
        RECT  5.430 1.065 5.505 1.155 ;
        RECT  5.340 0.505 5.430 1.155 ;
        RECT  5.310 1.265 5.410 1.515 ;
        RECT  5.210 0.505 5.340 0.615 ;
        RECT  4.570 0.905 5.340 0.995 ;
        RECT  4.960 1.265 5.310 1.355 ;
        RECT  4.300 0.705 5.240 0.815 ;
        RECT  4.780 1.085 5.180 1.175 ;
        RECT  5.030 0.305 5.120 0.585 ;
        RECT  4.690 0.495 5.030 0.585 ;
        RECT  4.870 1.265 4.960 1.525 ;
        RECT  4.055 1.435 4.870 1.525 ;
        RECT  4.680 1.085 4.780 1.310 ;
        RECT  4.600 0.305 4.690 0.585 ;
        RECT  4.480 1.200 4.680 1.310 ;
        RECT  4.180 0.305 4.600 0.415 ;
        RECT  4.435 0.905 4.570 1.090 ;
        RECT  4.185 0.525 4.300 1.325 ;
        RECT  4.050 0.525 4.185 0.640 ;
        RECT  3.940 0.905 4.080 1.035 ;
        RECT  3.965 1.255 4.055 1.525 ;
        RECT  2.575 1.255 3.965 1.345 ;
        RECT  3.700 0.275 3.960 0.385 ;
        RECT  3.830 0.520 3.940 1.165 ;
        RECT  3.700 1.435 3.875 1.545 ;
        RECT  3.525 0.520 3.830 0.630 ;
        RECT  3.625 1.045 3.830 1.165 ;
        RECT  3.535 0.740 3.740 0.870 ;
        RECT  0.690 0.275 3.700 0.365 ;
        RECT  1.955 1.435 3.700 1.525 ;
        RECT  3.445 0.740 3.535 1.165 ;
        RECT  3.150 1.045 3.445 1.165 ;
        RECT  3.040 0.455 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.675 2.755 1.165 ;
        RECT  2.665 0.490 2.670 1.165 ;
        RECT  2.560 0.490 2.665 0.765 ;
        RECT  2.485 0.890 2.575 1.345 ;
        RECT  2.055 0.675 2.560 0.765 ;
        RECT  2.170 0.890 2.485 1.000 ;
        RECT  1.210 0.475 2.435 0.585 ;
        RECT  2.280 1.130 2.395 1.305 ;
        RECT  1.600 1.215 2.280 1.305 ;
        RECT  1.945 0.675 2.055 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.945 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.245 1.215 1.600 1.345 ;
        RECT  1.330 1.015 1.520 1.125 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.905 0.510 0.910 0.835 ;
        RECT  0.795 0.510 0.905 1.345 ;
        RECT  0.720 0.510 0.795 0.620 ;
        RECT  0.400 1.000 0.795 1.090 ;
        RECT  0.475 0.265 0.690 0.365 ;
        RECT  0.535 1.250 0.645 1.525 ;
    END
END SEDFCNQD2

MACRO SEDFCNQD4
    CLASS CORE ;
    FOREIGN SEDFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.180 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0569 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.510 0.585 0.890 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.250 0.325 8.470 0.635 ;
        RECT  8.250 1.100 8.470 1.410 ;
        RECT  7.950 0.325 8.250 1.410 ;
        RECT  7.800 0.325 7.950 0.635 ;
        RECT  7.800 1.100 7.950 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0725 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.510 2.950 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.700 1.750 0.945 ;
        RECT  1.445 0.700 1.630 0.890 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.465 3.355 0.905 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.1094 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.710 7.150 0.890 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.710 -0.165 8.800 0.165 ;
        RECT  8.580 -0.165 8.710 0.670 ;
        RECT  7.710 -0.165 8.580 0.165 ;
        RECT  7.515 -0.165 7.710 0.420 ;
        RECT  6.625 -0.165 7.515 0.165 ;
        RECT  6.435 -0.165 6.625 0.400 ;
        RECT  4.995 -0.165 6.435 0.165 ;
        RECT  4.885 -0.165 4.995 0.405 ;
        RECT  0.185 -0.165 4.885 0.165 ;
        RECT  0.075 -0.165 0.185 0.465 ;
        RECT  0.000 -0.165 0.075 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.710 1.635 8.800 1.965 ;
        RECT  8.580 1.010 8.710 1.965 ;
        RECT  7.680 1.635 8.580 1.965 ;
        RECT  7.510 1.395 7.680 1.965 ;
        RECT  7.160 1.635 7.510 1.965 ;
        RECT  6.990 1.395 7.160 1.965 ;
        RECT  6.565 1.635 6.990 1.965 ;
        RECT  6.395 1.395 6.565 1.965 ;
        RECT  5.275 1.635 6.395 1.965 ;
        RECT  5.105 1.445 5.275 1.965 ;
        RECT  0.185 1.635 5.105 1.965 ;
        RECT  0.075 1.285 0.185 1.965 ;
        RECT  0.000 1.635 0.075 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.350 0.325 8.470 0.635 ;
        RECT  8.350 1.100 8.470 1.410 ;
        RECT  7.800 0.325 7.850 0.635 ;
        RECT  7.800 1.100 7.850 1.410 ;
        RECT  7.645 0.775 7.830 0.905 ;
        RECT  7.555 0.510 7.645 1.285 ;
        RECT  6.560 0.510 7.555 0.600 ;
        RECT  6.710 1.175 7.555 1.285 ;
        RECT  7.355 0.730 7.465 1.070 ;
        RECT  6.760 0.980 7.355 1.070 ;
        RECT  6.655 0.710 6.760 1.070 ;
        RECT  6.565 0.980 6.655 1.070 ;
        RECT  6.440 0.980 6.565 1.305 ;
        RECT  6.450 0.510 6.560 0.865 ;
        RECT  6.260 0.755 6.450 0.865 ;
        RECT  5.930 1.215 6.440 1.305 ;
        RECT  6.165 0.505 6.330 0.615 ;
        RECT  6.165 1.015 6.265 1.125 ;
        RECT  6.075 1.395 6.265 1.515 ;
        RECT  5.175 0.305 6.195 0.415 ;
        RECT  6.075 0.505 6.165 1.125 ;
        RECT  5.820 0.505 6.075 0.615 ;
        RECT  5.465 1.425 6.075 1.515 ;
        RECT  5.820 0.865 5.930 1.305 ;
        RECT  5.700 0.865 5.820 0.975 ;
        RECT  5.585 0.515 5.700 0.975 ;
        RECT  5.560 1.065 5.670 1.315 ;
        RECT  5.485 1.065 5.560 1.155 ;
        RECT  5.395 0.505 5.485 1.155 ;
        RECT  5.365 1.265 5.465 1.515 ;
        RECT  5.265 0.505 5.395 0.615 ;
        RECT  4.635 0.905 5.395 0.995 ;
        RECT  5.015 1.265 5.365 1.355 ;
        RECT  4.455 0.705 5.295 0.815 ;
        RECT  4.835 1.085 5.235 1.175 ;
        RECT  5.085 0.305 5.175 0.585 ;
        RECT  4.745 0.495 5.085 0.585 ;
        RECT  4.925 1.265 5.015 1.525 ;
        RECT  4.345 1.435 4.925 1.525 ;
        RECT  4.725 1.085 4.835 1.310 ;
        RECT  4.655 0.305 4.745 0.585 ;
        RECT  4.535 1.200 4.725 1.310 ;
        RECT  4.175 0.305 4.655 0.415 ;
        RECT  4.545 0.905 4.635 1.090 ;
        RECT  4.365 0.525 4.455 1.125 ;
        RECT  4.095 0.525 4.365 0.635 ;
        RECT  4.220 1.015 4.365 1.125 ;
        RECT  4.235 1.255 4.345 1.525 ;
        RECT  4.165 0.740 4.275 0.910 ;
        RECT  2.575 1.255 4.235 1.345 ;
        RECT  3.965 0.800 4.165 0.910 ;
        RECT  3.900 1.435 4.095 1.545 ;
        RECT  3.560 0.275 3.965 0.385 ;
        RECT  3.855 0.520 3.965 1.165 ;
        RECT  1.955 1.435 3.900 1.525 ;
        RECT  3.560 0.520 3.855 0.630 ;
        RECT  3.625 1.045 3.855 1.165 ;
        RECT  3.535 0.780 3.655 0.890 ;
        RECT  0.690 0.275 3.560 0.365 ;
        RECT  3.445 0.780 3.535 1.165 ;
        RECT  3.150 1.045 3.445 1.165 ;
        RECT  3.040 0.455 3.150 1.165 ;
        RECT  2.755 1.005 2.775 1.165 ;
        RECT  2.670 0.710 2.755 1.165 ;
        RECT  2.665 0.490 2.670 1.165 ;
        RECT  2.560 0.490 2.665 0.800 ;
        RECT  2.485 0.900 2.575 1.345 ;
        RECT  2.065 0.710 2.560 0.800 ;
        RECT  2.170 0.900 2.485 1.010 ;
        RECT  1.210 0.475 2.435 0.585 ;
        RECT  2.280 1.130 2.395 1.305 ;
        RECT  1.600 1.215 2.280 1.305 ;
        RECT  1.935 0.675 2.065 1.125 ;
        RECT  1.745 1.395 1.955 1.525 ;
        RECT  1.520 1.035 1.935 1.125 ;
        RECT  0.645 1.435 1.745 1.525 ;
        RECT  1.245 1.215 1.600 1.345 ;
        RECT  1.330 1.015 1.520 1.125 ;
        RECT  0.910 0.725 1.300 0.835 ;
        RECT  0.795 0.520 0.910 1.345 ;
        RECT  0.720 0.520 0.795 0.610 ;
        RECT  0.400 1.000 0.795 1.090 ;
        RECT  0.475 0.265 0.690 0.365 ;
        RECT  0.535 1.300 0.645 1.525 ;
    END
END SEDFCNQD4

MACRO SEDFD0
    CLASS CORE ;
    FOREIGN SEDFD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.485 6.950 1.290 ;
        RECT  6.815 0.485 6.850 0.665 ;
        RECT  6.815 1.040 6.850 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.080 6.435 1.190 ;
        RECT  6.350 0.475 6.405 0.685 ;
        RECT  6.250 0.475 6.350 1.190 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0495 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.815 -0.165 7.000 0.165 ;
        RECT  5.705 -0.165 5.815 0.385 ;
        RECT  2.110 -0.165 5.705 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 7.000 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.660 0.750 6.760 0.920 ;
        RECT  6.570 0.275 6.660 1.525 ;
        RECT  6.145 0.275 6.570 0.365 ;
        RECT  6.155 1.435 6.570 1.525 ;
        RECT  6.045 1.260 6.155 1.525 ;
        RECT  6.035 0.275 6.145 0.605 ;
        RECT  5.845 0.780 6.125 0.890 ;
        RECT  5.000 1.435 6.045 1.525 ;
        RECT  5.665 0.495 6.035 0.605 ;
        RECT  5.755 0.780 5.845 1.345 ;
        RECT  5.205 1.235 5.755 1.345 ;
        RECT  5.555 0.495 5.665 0.865 ;
        RECT  5.465 1.015 5.555 1.125 ;
        RECT  5.375 0.275 5.465 1.125 ;
        RECT  5.165 0.275 5.375 0.365 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.995 0.255 5.165 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.995 0.365 ;
        RECT  4.890 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.800 0.735 4.845 0.905 ;
        RECT  4.710 0.475 4.800 0.905 ;
        RECT  4.365 0.475 4.710 0.565 ;
        RECT  4.505 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.740 3.655 0.910 ;
        RECT  3.440 0.515 3.530 1.165 ;
        RECT  3.135 0.515 3.440 0.620 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.305 0.360 1.090 ;
        RECT  0.045 0.305 0.270 0.415 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFD0

MACRO SEDFD1
    CLASS CORE ;
    FOREIGN SEDFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.285 6.950 1.490 ;
        RECT  6.815 0.285 6.850 0.665 ;
        RECT  6.815 1.050 6.850 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.080 6.435 1.190 ;
        RECT  6.350 0.475 6.405 0.685 ;
        RECT  6.250 0.475 6.350 1.190 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.815 -0.165 7.000 0.165 ;
        RECT  5.705 -0.165 5.815 0.385 ;
        RECT  2.110 -0.165 5.705 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 7.000 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.660 0.750 6.760 0.920 ;
        RECT  6.570 0.275 6.660 1.525 ;
        RECT  6.160 0.275 6.570 0.365 ;
        RECT  6.155 1.435 6.570 1.525 ;
        RECT  6.050 0.275 6.160 0.605 ;
        RECT  6.045 1.260 6.155 1.525 ;
        RECT  5.845 0.780 6.125 0.890 ;
        RECT  5.665 0.495 6.050 0.605 ;
        RECT  5.000 1.435 6.045 1.525 ;
        RECT  5.755 0.780 5.845 1.345 ;
        RECT  5.205 1.235 5.755 1.345 ;
        RECT  5.555 0.495 5.665 0.865 ;
        RECT  5.465 1.015 5.555 1.125 ;
        RECT  5.375 0.275 5.465 1.125 ;
        RECT  5.165 0.275 5.375 0.365 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.995 0.255 5.165 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.995 0.365 ;
        RECT  4.890 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.800 0.735 4.845 0.905 ;
        RECT  4.710 0.475 4.800 0.905 ;
        RECT  4.365 0.475 4.710 0.565 ;
        RECT  4.505 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.225 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.740 3.655 0.910 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFD1

MACRO SEDFD2
    CLASS CORE ;
    FOREIGN SEDFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.285 7.150 1.490 ;
        RECT  6.965 0.285 7.050 0.665 ;
        RECT  6.965 1.050 7.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.550 0.475 6.575 0.685 ;
        RECT  6.550 1.155 6.575 1.325 ;
        RECT  6.450 0.475 6.550 1.325 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.775 -0.165 7.400 0.165 ;
        RECT  5.665 -0.165 5.775 0.385 ;
        RECT  2.110 -0.165 5.665 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 7.400 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.810 0.750 6.920 0.920 ;
        RECT  6.720 0.275 6.810 1.525 ;
        RECT  6.100 0.275 6.720 0.365 ;
        RECT  6.100 1.435 6.720 1.525 ;
        RECT  5.845 0.780 6.330 0.890 ;
        RECT  5.990 0.275 6.100 0.605 ;
        RECT  5.990 1.150 6.100 1.525 ;
        RECT  5.665 0.495 5.990 0.605 ;
        RECT  5.000 1.435 5.990 1.525 ;
        RECT  5.755 0.780 5.845 1.345 ;
        RECT  5.205 1.235 5.755 1.345 ;
        RECT  5.555 0.495 5.665 0.865 ;
        RECT  5.465 1.015 5.555 1.125 ;
        RECT  5.375 0.275 5.465 1.125 ;
        RECT  5.165 0.275 5.375 0.365 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.995 0.255 5.165 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.995 0.365 ;
        RECT  4.890 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.800 0.735 4.845 0.905 ;
        RECT  4.710 0.475 4.800 0.905 ;
        RECT  4.365 0.475 4.710 0.565 ;
        RECT  4.505 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.740 3.655 0.910 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFD2

MACRO SEDFD4
    CLASS CORE ;
    FOREIGN SEDFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.450 0.325 8.705 0.635 ;
        RECT  8.450 1.100 8.705 1.410 ;
        RECT  8.150 0.325 8.450 1.410 ;
        RECT  8.035 0.325 8.150 0.635 ;
        RECT  8.035 1.100 8.150 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.515 7.705 0.685 ;
        RECT  7.450 1.115 7.705 1.285 ;
        RECT  7.150 0.515 7.450 1.285 ;
        RECT  7.035 0.515 7.150 0.685 ;
        RECT  7.035 1.115 7.150 1.285 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.375 -0.165 9.000 0.165 ;
        RECT  6.265 -0.165 6.375 0.385 ;
        RECT  2.110 -0.165 6.265 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.330 1.635 9.000 1.965 ;
        RECT  5.160 1.445 5.330 1.965 ;
        RECT  4.760 1.635 5.160 1.965 ;
        RECT  4.590 1.445 4.760 1.965 ;
        RECT  0.525 1.635 4.590 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.550 0.325 8.705 0.635 ;
        RECT  8.550 1.100 8.705 1.410 ;
        RECT  8.035 0.325 8.050 0.635 ;
        RECT  8.035 1.100 8.050 1.410 ;
        RECT  7.550 0.515 7.705 0.685 ;
        RECT  7.550 1.115 7.705 1.285 ;
        RECT  7.035 0.515 7.050 0.685 ;
        RECT  7.035 1.115 7.050 1.285 ;
        RECT  7.910 0.750 8.020 0.920 ;
        RECT  7.820 0.275 7.910 1.525 ;
        RECT  6.695 0.275 7.820 0.365 ;
        RECT  6.700 1.435 7.820 1.525 ;
        RECT  6.445 0.780 6.930 0.890 ;
        RECT  6.590 1.060 6.700 1.525 ;
        RECT  6.585 0.275 6.695 0.670 ;
        RECT  5.590 1.435 6.590 1.525 ;
        RECT  6.265 0.560 6.585 0.670 ;
        RECT  6.355 0.780 6.445 1.345 ;
        RECT  5.865 1.235 6.355 1.345 ;
        RECT  6.155 0.560 6.265 0.865 ;
        RECT  6.065 1.015 6.155 1.125 ;
        RECT  5.975 0.275 6.065 1.125 ;
        RECT  5.765 0.275 5.975 0.365 ;
        RECT  5.865 0.465 5.885 0.575 ;
        RECT  5.755 0.465 5.865 1.345 ;
        RECT  5.595 0.255 5.765 0.365 ;
        RECT  5.715 0.465 5.755 0.575 ;
        RECT  5.590 1.065 5.635 1.175 ;
        RECT  4.435 0.275 5.595 0.365 ;
        RECT  5.450 0.455 5.590 1.175 ;
        RECT  5.500 1.265 5.590 1.525 ;
        RECT  4.340 1.265 5.500 1.355 ;
        RECT  5.010 0.455 5.450 0.555 ;
        RECT  4.615 1.065 5.450 1.175 ;
        RECT  4.795 0.765 5.030 0.875 ;
        RECT  4.910 0.455 5.010 0.645 ;
        RECT  4.705 0.475 4.795 0.875 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.175 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.750 3.655 0.920 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.305 0.360 1.090 ;
        RECT  0.045 0.305 0.270 0.415 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFD4

MACRO SEDFKCND0
    CLASS CORE ;
    FOREIGN SEDFKCND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0189 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.900 2.760 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0528 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.445 0.910 3.750 1.090 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.475 7.750 1.290 ;
        RECT  7.620 0.475 7.650 0.675 ;
        RECT  7.620 1.020 7.650 1.290 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.490 7.350 1.230 ;
        RECT  7.125 0.490 7.250 0.660 ;
        RECT  7.125 1.020 7.250 1.230 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0439 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.190 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0428 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.810 1.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0227 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.900 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.385 -0.165 7.800 0.165 ;
        RECT  5.385 0.475 5.555 0.585 ;
        RECT  5.285 -0.165 5.385 0.585 ;
        RECT  2.865 -0.165 5.285 0.165 ;
        RECT  2.760 -0.165 2.865 0.590 ;
        RECT  0.000 -0.165 2.760 0.165 ;
        RECT  2.535 0.480 2.760 0.590 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.470 1.635 7.800 1.965 ;
        RECT  7.300 1.515 7.470 1.965 ;
        RECT  5.590 1.635 7.300 1.965 ;
        RECT  5.400 1.435 5.590 1.965 ;
        RECT  2.820 1.635 5.400 1.965 ;
        RECT  2.675 1.385 2.820 1.965 ;
        RECT  0.445 1.635 2.675 1.965 ;
        RECT  0.335 1.250 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.530 0.755 7.560 0.925 ;
        RECT  7.440 0.285 7.530 1.425 ;
        RECT  6.410 0.285 7.440 0.385 ;
        RECT  6.955 1.335 7.440 1.425 ;
        RECT  7.015 0.785 7.100 0.895 ;
        RECT  6.925 0.505 7.015 1.230 ;
        RECT  6.855 1.335 6.955 1.495 ;
        RECT  6.565 0.505 6.925 0.615 ;
        RECT  6.835 1.110 6.925 1.230 ;
        RECT  5.850 1.395 6.855 1.495 ;
        RECT  6.745 0.755 6.820 0.925 ;
        RECT  6.655 0.755 6.745 1.305 ;
        RECT  6.085 1.215 6.655 1.305 ;
        RECT  6.455 0.505 6.565 1.120 ;
        RECT  6.295 0.255 6.410 0.425 ;
        RECT  6.205 0.585 6.315 1.120 ;
        RECT  6.115 0.275 6.205 0.675 ;
        RECT  5.975 0.275 6.115 0.365 ;
        RECT  6.025 0.830 6.085 1.305 ;
        RECT  5.980 0.505 6.025 1.305 ;
        RECT  5.915 0.505 5.980 0.930 ;
        RECT  5.770 0.255 5.975 0.365 ;
        RECT  5.820 1.020 5.890 1.140 ;
        RECT  5.740 1.230 5.850 1.495 ;
        RECT  5.765 0.675 5.820 1.140 ;
        RECT  5.720 0.465 5.765 1.140 ;
        RECT  5.265 1.230 5.740 1.330 ;
        RECT  5.655 0.465 5.720 0.765 ;
        RECT  5.380 0.675 5.655 0.765 ;
        RECT  5.520 0.875 5.630 1.120 ;
        RECT  5.065 1.030 5.520 1.120 ;
        RECT  5.260 0.675 5.380 0.915 ;
        RECT  5.175 1.230 5.265 1.525 ;
        RECT  3.040 1.435 5.175 1.525 ;
        RECT  5.020 1.030 5.065 1.345 ;
        RECT  4.955 0.300 5.020 1.345 ;
        RECT  4.910 0.300 4.955 1.120 ;
        RECT  4.665 1.215 4.850 1.345 ;
        RECT  4.670 0.520 4.785 1.125 ;
        RECT  4.595 0.255 4.765 0.365 ;
        RECT  4.420 0.520 4.670 0.635 ;
        RECT  4.420 1.015 4.670 1.125 ;
        RECT  3.335 1.255 4.665 1.345 ;
        RECT  3.290 0.275 4.595 0.365 ;
        RECT  4.330 0.775 4.445 0.895 ;
        RECT  4.240 0.500 4.330 1.145 ;
        RECT  3.860 0.500 4.240 0.610 ;
        RECT  3.875 1.035 4.240 1.145 ;
        RECT  3.510 0.600 3.640 0.790 ;
        RECT  3.210 0.700 3.510 0.790 ;
        RECT  3.130 1.215 3.335 1.345 ;
        RECT  3.160 0.275 3.290 0.560 ;
        RECT  3.040 0.700 3.210 1.090 ;
        RECT  2.445 0.700 3.040 0.790 ;
        RECT  2.940 1.205 3.040 1.525 ;
        RECT  2.585 1.205 2.940 1.295 ;
        RECT  2.495 1.205 2.585 1.525 ;
        RECT  1.450 1.435 2.495 1.525 ;
        RECT  2.350 0.480 2.445 0.790 ;
        RECT  2.350 1.175 2.405 1.345 ;
        RECT  2.260 0.480 2.350 1.345 ;
        RECT  2.170 0.265 2.290 0.375 ;
        RECT  2.080 0.265 2.170 1.340 ;
        RECT  2.050 0.265 2.080 0.655 ;
        RECT  2.030 1.170 2.080 1.340 ;
        RECT  1.960 0.750 1.990 0.920 ;
        RECT  1.850 0.495 1.960 1.080 ;
        RECT  1.265 0.495 1.850 0.600 ;
        RECT  1.655 0.990 1.850 1.080 ;
        RECT  1.495 0.275 1.705 0.405 ;
        RECT  1.545 0.990 1.655 1.345 ;
        RECT  0.725 0.275 1.495 0.365 ;
        RECT  1.360 1.010 1.450 1.525 ;
        RECT  1.175 0.475 1.265 1.330 ;
        RECT  1.095 0.475 1.175 0.665 ;
        RECT  0.955 1.240 1.175 1.330 ;
        RECT  0.990 0.875 1.085 1.085 ;
        RECT  0.900 0.525 0.990 1.085 ;
        RECT  0.845 1.240 0.955 1.515 ;
        RECT  0.540 0.525 0.900 0.615 ;
        RECT  0.555 0.275 0.725 0.415 ;
        RECT  0.435 0.525 0.540 1.140 ;
        RECT  0.410 0.325 0.435 1.140 ;
        RECT  0.325 0.325 0.410 0.625 ;
        RECT  0.185 1.040 0.410 1.140 ;
        RECT  0.075 1.040 0.185 1.430 ;
    END
END SEDFKCND0

MACRO SEDFKCND1
    CLASS CORE ;
    FOREIGN SEDFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.900 2.760 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0580 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.800 3.495 1.120 ;
        RECT  3.350 0.800 3.385 0.890 ;
        RECT  3.045 0.710 3.350 0.890 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 0.275 7.950 1.490 ;
        RECT  7.820 0.275 7.850 0.675 ;
        RECT  7.820 1.020 7.850 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1510 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.490 7.550 1.230 ;
        RECT  7.325 0.490 7.450 0.660 ;
        RECT  7.325 1.020 7.450 1.230 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.190 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.810 1.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.900 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.585 -0.165 8.000 0.165 ;
        RECT  5.585 0.475 5.755 0.585 ;
        RECT  5.485 -0.165 5.585 0.585 ;
        RECT  2.865 -0.165 5.485 0.165 ;
        RECT  2.760 -0.165 2.865 0.600 ;
        RECT  0.000 -0.165 2.760 0.165 ;
        RECT  2.525 0.490 2.760 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.790 1.635 8.000 1.965 ;
        RECT  5.600 1.435 5.790 1.965 ;
        RECT  2.820 1.635 5.600 1.965 ;
        RECT  2.675 1.385 2.820 1.965 ;
        RECT  0.445 1.635 2.675 1.965 ;
        RECT  0.335 1.250 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.730 0.755 7.760 0.925 ;
        RECT  7.640 0.285 7.730 1.435 ;
        RECT  6.610 0.285 7.640 0.385 ;
        RECT  7.155 1.335 7.640 1.435 ;
        RECT  7.215 0.785 7.300 0.895 ;
        RECT  7.125 0.505 7.215 1.230 ;
        RECT  7.055 1.335 7.155 1.495 ;
        RECT  6.765 0.505 7.125 0.615 ;
        RECT  7.035 1.110 7.125 1.230 ;
        RECT  6.050 1.395 7.055 1.495 ;
        RECT  6.945 0.755 7.020 0.925 ;
        RECT  6.855 0.755 6.945 1.305 ;
        RECT  6.285 1.215 6.855 1.305 ;
        RECT  6.655 0.505 6.765 1.120 ;
        RECT  6.495 0.255 6.610 0.425 ;
        RECT  6.405 0.585 6.515 1.120 ;
        RECT  6.315 0.275 6.405 0.675 ;
        RECT  6.175 0.275 6.315 0.365 ;
        RECT  6.225 0.830 6.285 1.305 ;
        RECT  6.180 0.505 6.225 1.305 ;
        RECT  6.115 0.505 6.180 0.930 ;
        RECT  5.970 0.255 6.175 0.365 ;
        RECT  6.020 1.020 6.090 1.140 ;
        RECT  5.940 1.230 6.050 1.495 ;
        RECT  5.965 0.675 6.020 1.140 ;
        RECT  5.920 0.465 5.965 1.140 ;
        RECT  5.465 1.230 5.940 1.330 ;
        RECT  5.855 0.465 5.920 0.765 ;
        RECT  5.580 0.675 5.855 0.765 ;
        RECT  5.720 0.875 5.830 1.120 ;
        RECT  5.265 1.030 5.720 1.120 ;
        RECT  5.460 0.675 5.580 0.915 ;
        RECT  5.375 1.230 5.465 1.525 ;
        RECT  3.040 1.435 5.375 1.525 ;
        RECT  5.220 1.030 5.265 1.345 ;
        RECT  5.155 0.300 5.220 1.345 ;
        RECT  5.110 0.300 5.155 1.120 ;
        RECT  4.865 1.215 5.050 1.345 ;
        RECT  4.870 0.520 4.985 1.125 ;
        RECT  4.795 0.255 4.965 0.365 ;
        RECT  4.560 0.520 4.870 0.635 ;
        RECT  4.620 1.015 4.870 1.125 ;
        RECT  3.395 1.255 4.865 1.345 ;
        RECT  3.310 0.275 4.795 0.365 ;
        RECT  4.350 0.775 4.645 0.895 ;
        RECT  4.260 0.500 4.350 1.145 ;
        RECT  4.000 0.500 4.260 0.610 ;
        RECT  4.075 1.035 4.260 1.145 ;
        RECT  3.615 0.600 3.725 1.165 ;
        RECT  3.555 0.600 3.615 0.690 ;
        RECT  3.445 0.475 3.555 0.690 ;
        RECT  3.190 1.215 3.395 1.345 ;
        RECT  3.140 0.275 3.310 0.585 ;
        RECT  2.940 0.990 3.240 1.090 ;
        RECT  2.940 1.205 3.040 1.525 ;
        RECT  2.850 0.700 2.940 1.090 ;
        RECT  2.585 1.205 2.940 1.295 ;
        RECT  2.435 0.700 2.850 0.790 ;
        RECT  2.495 1.205 2.585 1.525 ;
        RECT  1.450 1.435 2.495 1.525 ;
        RECT  2.350 0.475 2.435 0.790 ;
        RECT  2.350 1.175 2.405 1.345 ;
        RECT  2.260 0.475 2.350 1.345 ;
        RECT  2.170 0.265 2.290 0.375 ;
        RECT  2.080 0.265 2.170 1.340 ;
        RECT  2.050 0.265 2.080 0.655 ;
        RECT  2.030 1.170 2.080 1.340 ;
        RECT  1.960 0.750 1.990 0.920 ;
        RECT  1.850 0.495 1.960 1.080 ;
        RECT  1.265 0.495 1.850 0.600 ;
        RECT  1.655 0.990 1.850 1.080 ;
        RECT  1.495 0.275 1.705 0.405 ;
        RECT  1.545 0.990 1.655 1.345 ;
        RECT  0.735 0.275 1.495 0.365 ;
        RECT  1.360 1.010 1.450 1.525 ;
        RECT  1.175 0.475 1.265 1.330 ;
        RECT  1.095 0.475 1.175 0.665 ;
        RECT  0.955 1.240 1.175 1.330 ;
        RECT  0.990 0.875 1.085 1.085 ;
        RECT  0.900 0.525 0.990 1.085 ;
        RECT  0.845 1.240 0.955 1.515 ;
        RECT  0.530 0.525 0.900 0.615 ;
        RECT  0.555 0.275 0.735 0.405 ;
        RECT  0.435 0.525 0.530 1.140 ;
        RECT  0.420 0.315 0.435 1.140 ;
        RECT  0.325 0.315 0.420 0.625 ;
        RECT  0.185 1.040 0.420 1.140 ;
        RECT  0.075 1.040 0.185 1.420 ;
    END
END SEDFKCND1

MACRO SEDFKCND2
    CLASS CORE ;
    FOREIGN SEDFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0203 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.900 2.760 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0580 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.800 3.495 1.120 ;
        RECT  3.350 0.800 3.385 0.890 ;
        RECT  3.045 0.710 3.350 0.890 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 0.275 8.150 1.490 ;
        RECT  7.965 0.275 8.050 0.675 ;
        RECT  7.965 1.020 8.050 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.550 0.490 7.575 0.680 ;
        RECT  7.550 1.080 7.575 1.290 ;
        RECT  7.450 0.490 7.550 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.190 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.810 1.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.900 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.525 -0.165 8.400 0.165 ;
        RECT  5.525 0.475 5.695 0.585 ;
        RECT  5.425 -0.165 5.525 0.585 ;
        RECT  2.865 -0.165 5.425 0.165 ;
        RECT  2.760 -0.165 2.865 0.600 ;
        RECT  0.000 -0.165 2.760 0.165 ;
        RECT  2.525 0.490 2.760 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 1.635 8.400 1.965 ;
        RECT  5.540 1.435 5.730 1.965 ;
        RECT  2.820 1.635 5.540 1.965 ;
        RECT  2.675 1.385 2.820 1.965 ;
        RECT  0.445 1.635 2.675 1.965 ;
        RECT  0.335 1.250 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.875 0.755 7.910 0.925 ;
        RECT  7.785 0.285 7.875 1.495 ;
        RECT  6.550 0.285 7.785 0.385 ;
        RECT  5.990 1.395 7.785 1.495 ;
        RECT  7.155 0.785 7.340 0.895 ;
        RECT  7.065 0.505 7.155 1.305 ;
        RECT  6.705 0.505 7.065 0.615 ;
        RECT  6.985 1.115 7.065 1.305 ;
        RECT  6.885 0.755 6.960 0.925 ;
        RECT  6.795 0.755 6.885 1.305 ;
        RECT  6.225 1.215 6.795 1.305 ;
        RECT  6.595 0.505 6.705 1.120 ;
        RECT  6.435 0.255 6.550 0.425 ;
        RECT  6.345 0.585 6.455 1.120 ;
        RECT  6.255 0.275 6.345 0.675 ;
        RECT  6.115 0.275 6.255 0.365 ;
        RECT  6.165 0.830 6.225 1.305 ;
        RECT  6.120 0.505 6.165 1.305 ;
        RECT  6.055 0.505 6.120 0.930 ;
        RECT  5.910 0.255 6.115 0.365 ;
        RECT  5.960 1.020 6.030 1.140 ;
        RECT  5.880 1.230 5.990 1.495 ;
        RECT  5.905 0.675 5.960 1.140 ;
        RECT  5.860 0.465 5.905 1.140 ;
        RECT  5.405 1.230 5.880 1.330 ;
        RECT  5.795 0.465 5.860 0.765 ;
        RECT  5.520 0.675 5.795 0.765 ;
        RECT  5.660 0.875 5.770 1.120 ;
        RECT  5.205 1.030 5.660 1.120 ;
        RECT  5.400 0.675 5.520 0.915 ;
        RECT  5.315 1.230 5.405 1.525 ;
        RECT  3.040 1.435 5.315 1.525 ;
        RECT  5.160 1.030 5.205 1.345 ;
        RECT  5.095 0.300 5.160 1.345 ;
        RECT  5.050 0.300 5.095 1.120 ;
        RECT  4.805 1.215 4.990 1.345 ;
        RECT  4.810 0.520 4.925 1.125 ;
        RECT  4.735 0.255 4.905 0.365 ;
        RECT  4.500 0.520 4.810 0.635 ;
        RECT  4.580 1.015 4.810 1.125 ;
        RECT  3.395 1.255 4.805 1.345 ;
        RECT  3.310 0.275 4.735 0.365 ;
        RECT  4.350 0.775 4.590 0.895 ;
        RECT  4.260 0.500 4.350 1.145 ;
        RECT  4.000 0.500 4.260 0.610 ;
        RECT  4.070 1.035 4.260 1.145 ;
        RECT  3.615 0.600 3.725 1.165 ;
        RECT  3.555 0.600 3.615 0.690 ;
        RECT  3.445 0.475 3.555 0.690 ;
        RECT  3.190 1.215 3.395 1.345 ;
        RECT  3.140 0.275 3.310 0.585 ;
        RECT  2.940 0.990 3.240 1.090 ;
        RECT  2.940 1.205 3.040 1.525 ;
        RECT  2.850 0.700 2.940 1.090 ;
        RECT  2.585 1.205 2.940 1.295 ;
        RECT  2.435 0.700 2.850 0.790 ;
        RECT  2.495 1.205 2.585 1.525 ;
        RECT  1.450 1.435 2.495 1.525 ;
        RECT  2.350 0.475 2.435 0.790 ;
        RECT  2.350 1.175 2.405 1.345 ;
        RECT  2.260 0.475 2.350 1.345 ;
        RECT  2.170 0.265 2.290 0.375 ;
        RECT  2.080 0.265 2.170 1.340 ;
        RECT  2.050 0.265 2.080 0.655 ;
        RECT  2.030 1.170 2.080 1.340 ;
        RECT  1.960 0.750 1.990 0.920 ;
        RECT  1.850 0.495 1.960 1.080 ;
        RECT  1.265 0.495 1.850 0.600 ;
        RECT  1.655 0.990 1.850 1.080 ;
        RECT  1.495 0.275 1.705 0.405 ;
        RECT  1.545 0.990 1.655 1.345 ;
        RECT  0.725 0.275 1.495 0.365 ;
        RECT  1.360 1.010 1.450 1.525 ;
        RECT  1.175 0.475 1.265 1.330 ;
        RECT  1.095 0.475 1.175 0.665 ;
        RECT  0.955 1.240 1.175 1.330 ;
        RECT  0.990 0.875 1.085 1.085 ;
        RECT  0.900 0.525 0.990 1.085 ;
        RECT  0.845 1.240 0.955 1.515 ;
        RECT  0.530 0.525 0.900 0.615 ;
        RECT  0.555 0.275 0.725 0.405 ;
        RECT  0.435 0.525 0.530 1.140 ;
        RECT  0.420 0.315 0.435 1.140 ;
        RECT  0.325 0.315 0.420 0.625 ;
        RECT  0.185 1.040 0.420 1.140 ;
        RECT  0.075 1.040 0.185 1.420 ;
    END
END SEDFKCND2

MACRO SEDFKCND4
    CLASS CORE ;
    FOREIGN SEDFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.900 2.760 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0581 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 0.800 3.450 1.120 ;
        RECT  3.340 0.710 3.350 1.120 ;
        RECT  3.045 0.710 3.340 0.890 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.250 0.325 9.505 0.635 ;
        RECT  9.250 1.100 9.505 1.410 ;
        RECT  8.950 0.325 9.250 1.410 ;
        RECT  8.835 0.325 8.950 0.635 ;
        RECT  8.835 1.100 8.950 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.250 0.485 8.505 0.655 ;
        RECT  8.250 1.070 8.505 1.240 ;
        RECT  7.950 0.485 8.250 1.240 ;
        RECT  7.815 0.485 7.950 0.655 ;
        RECT  7.815 1.070 7.950 1.240 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.190 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.810 1.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.900 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.480 -0.165 9.800 0.165 ;
        RECT  5.480 0.475 5.650 0.585 ;
        RECT  5.380 -0.165 5.480 0.585 ;
        RECT  2.865 -0.165 5.380 0.165 ;
        RECT  2.760 -0.165 2.865 0.600 ;
        RECT  0.000 -0.165 2.760 0.165 ;
        RECT  2.510 0.490 2.760 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 1.635 9.800 1.965 ;
        RECT  5.495 1.435 5.685 1.965 ;
        RECT  2.820 1.635 5.495 1.965 ;
        RECT  2.675 1.385 2.820 1.965 ;
        RECT  0.445 1.635 2.675 1.965 ;
        RECT  0.335 1.250 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.350 0.325 9.505 0.635 ;
        RECT  9.350 1.100 9.505 1.410 ;
        RECT  8.835 0.325 8.850 0.635 ;
        RECT  8.835 1.100 8.850 1.410 ;
        RECT  8.350 0.485 8.505 0.655 ;
        RECT  8.350 1.070 8.505 1.240 ;
        RECT  7.815 0.485 7.850 0.655 ;
        RECT  7.815 1.070 7.850 1.240 ;
        RECT  8.730 0.750 8.810 0.920 ;
        RECT  8.620 0.285 8.730 1.495 ;
        RECT  6.985 0.285 8.620 0.375 ;
        RECT  6.985 1.385 8.620 1.495 ;
        RECT  7.710 0.750 7.820 0.920 ;
        RECT  7.705 0.485 7.710 0.920 ;
        RECT  7.605 0.485 7.705 1.265 ;
        RECT  7.210 0.485 7.605 0.610 ;
        RECT  7.315 1.155 7.605 1.265 ;
        RECT  7.365 0.745 7.475 1.045 ;
        RECT  6.240 0.955 7.365 1.045 ;
        RECT  7.120 0.485 7.210 0.865 ;
        RECT  6.825 0.765 7.120 0.865 ;
        RECT  6.855 0.285 6.985 0.665 ;
        RECT  6.855 1.145 6.985 1.495 ;
        RECT  6.380 0.285 6.855 0.375 ;
        RECT  6.530 1.395 6.855 1.495 ;
        RECT  6.360 1.135 6.530 1.495 ;
        RECT  6.270 0.285 6.380 0.705 ;
        RECT  5.945 1.395 6.360 1.495 ;
        RECT  6.130 0.830 6.240 1.265 ;
        RECT  6.120 0.830 6.130 0.930 ;
        RECT  6.010 0.505 6.120 0.930 ;
        RECT  5.915 1.060 5.985 1.165 ;
        RECT  5.835 1.255 5.945 1.495 ;
        RECT  5.860 0.675 5.915 1.165 ;
        RECT  5.815 0.465 5.860 1.165 ;
        RECT  5.360 1.255 5.835 1.345 ;
        RECT  5.750 0.465 5.815 0.765 ;
        RECT  5.475 0.675 5.750 0.765 ;
        RECT  5.615 0.875 5.725 1.120 ;
        RECT  5.160 1.030 5.615 1.120 ;
        RECT  5.355 0.675 5.475 0.915 ;
        RECT  5.270 1.255 5.360 1.525 ;
        RECT  3.040 1.435 5.270 1.525 ;
        RECT  5.115 1.030 5.160 1.345 ;
        RECT  5.050 0.300 5.115 1.345 ;
        RECT  5.005 0.300 5.050 1.120 ;
        RECT  4.760 1.215 4.945 1.345 ;
        RECT  4.765 0.520 4.880 1.125 ;
        RECT  4.690 0.255 4.860 0.365 ;
        RECT  4.455 0.520 4.765 0.635 ;
        RECT  4.535 1.015 4.765 1.125 ;
        RECT  3.395 1.255 4.760 1.345 ;
        RECT  3.310 0.275 4.690 0.365 ;
        RECT  4.350 0.775 4.545 0.895 ;
        RECT  4.260 0.500 4.350 1.145 ;
        RECT  3.955 0.500 4.260 0.610 ;
        RECT  4.030 1.035 4.260 1.145 ;
        RECT  3.570 0.600 3.680 1.165 ;
        RECT  3.555 0.600 3.570 0.690 ;
        RECT  3.445 0.475 3.555 0.690 ;
        RECT  3.190 1.215 3.395 1.345 ;
        RECT  3.140 0.275 3.310 0.585 ;
        RECT  2.940 0.980 3.240 1.090 ;
        RECT  2.940 1.205 3.040 1.525 ;
        RECT  2.850 0.700 2.940 1.090 ;
        RECT  2.585 1.205 2.940 1.295 ;
        RECT  2.390 0.700 2.850 0.790 ;
        RECT  2.495 1.205 2.585 1.525 ;
        RECT  1.450 1.435 2.495 1.525 ;
        RECT  2.350 1.175 2.405 1.345 ;
        RECT  2.350 0.475 2.390 0.790 ;
        RECT  2.260 0.475 2.350 1.345 ;
        RECT  2.170 0.265 2.275 0.375 ;
        RECT  2.080 0.265 2.170 1.340 ;
        RECT  2.030 0.265 2.080 0.655 ;
        RECT  2.030 1.170 2.080 1.340 ;
        RECT  1.940 0.750 1.990 0.920 ;
        RECT  1.850 0.495 1.940 1.080 ;
        RECT  1.265 0.495 1.850 0.600 ;
        RECT  1.655 0.990 1.850 1.080 ;
        RECT  1.480 0.275 1.690 0.405 ;
        RECT  1.545 0.990 1.655 1.345 ;
        RECT  0.725 0.275 1.480 0.365 ;
        RECT  1.360 1.010 1.450 1.525 ;
        RECT  1.175 0.475 1.265 1.330 ;
        RECT  1.080 0.475 1.175 0.665 ;
        RECT  0.955 1.240 1.175 1.330 ;
        RECT  0.990 0.875 1.085 1.085 ;
        RECT  0.900 0.525 0.990 1.085 ;
        RECT  0.845 1.240 0.955 1.515 ;
        RECT  0.530 0.525 0.900 0.615 ;
        RECT  0.555 0.275 0.725 0.405 ;
        RECT  0.435 0.525 0.530 1.140 ;
        RECT  0.420 0.315 0.435 1.140 ;
        RECT  0.325 0.315 0.420 0.625 ;
        RECT  0.185 1.040 0.420 1.140 ;
        RECT  0.075 1.040 0.185 1.420 ;
    END
END SEDFKCND4

MACRO SEDFKCNQD0
    CLASS CORE ;
    FOREIGN SEDFKCNQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.445 0.710 3.755 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0561 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.955 0.510 2.010 0.815 ;
        RECT  1.900 0.510 1.955 1.090 ;
        RECT  1.845 0.710 1.900 1.090 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0399 ;
        ANTENNADIFFAREA 0.1430 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.275 6.950 1.525 ;
        RECT  6.815 0.275 6.850 0.650 ;
        RECT  6.815 1.055 6.850 1.525 ;
        RECT  6.485 0.560 6.815 0.650 ;
        RECT  5.855 1.435 6.815 1.525 ;
        RECT  6.375 0.560 6.485 0.905 ;
        RECT  5.765 1.265 5.855 1.525 ;
        RECT  5.295 1.265 5.765 1.355 ;
        RECT  5.205 1.265 5.295 1.525 ;
        RECT  1.465 1.435 5.205 1.525 ;
        RECT  1.355 0.990 1.465 1.525 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0414 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.355 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0273 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.785 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.845 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.510 1.750 0.700 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.600 -0.165 7.000 0.165 ;
        RECT  6.490 -0.165 6.600 0.450 ;
        RECT  2.515 -0.165 6.490 0.165 ;
        RECT  2.375 -0.165 2.515 0.605 ;
        RECT  0.000 -0.165 2.375 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.595 1.635 7.000 1.965 ;
        RECT  5.425 1.445 5.595 1.965 ;
        RECT  0.475 1.635 5.425 1.965 ;
        RECT  0.305 1.200 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.715 0.750 6.760 0.920 ;
        RECT  6.615 0.750 6.715 1.345 ;
        RECT  6.075 1.235 6.615 1.345 ;
        RECT  6.255 1.025 6.395 1.135 ;
        RECT  6.165 0.275 6.255 1.135 ;
        RECT  6.030 0.275 6.165 0.365 ;
        RECT  5.975 0.475 6.075 1.345 ;
        RECT  5.820 0.255 6.030 0.365 ;
        RECT  5.765 0.505 5.875 1.175 ;
        RECT  5.245 0.275 5.820 0.365 ;
        RECT  5.445 0.505 5.765 0.620 ;
        RECT  5.650 0.740 5.675 0.910 ;
        RECT  5.560 0.740 5.650 1.175 ;
        RECT  5.065 1.085 5.560 1.175 ;
        RECT  5.335 0.505 5.445 0.940 ;
        RECT  5.035 0.255 5.245 0.365 ;
        RECT  5.050 0.485 5.065 1.175 ;
        RECT  4.940 0.485 5.050 1.270 ;
        RECT  4.530 0.795 4.820 0.925 ;
        RECT  4.680 0.275 4.790 0.480 ;
        RECT  4.680 1.070 4.790 1.345 ;
        RECT  2.970 0.275 4.680 0.365 ;
        RECT  2.740 1.255 4.680 1.345 ;
        RECT  4.420 0.475 4.530 1.165 ;
        RECT  4.240 0.490 4.330 1.165 ;
        RECT  3.840 0.490 4.240 0.600 ;
        RECT  3.840 1.065 4.240 1.165 ;
        RECT  3.305 0.490 3.730 0.600 ;
        RECT  3.305 1.065 3.730 1.165 ;
        RECT  3.195 0.490 3.305 1.165 ;
        RECT  2.935 0.725 3.045 1.090 ;
        RECT  2.840 0.275 2.970 0.605 ;
        RECT  2.260 0.725 2.935 0.815 ;
        RECT  2.605 0.925 2.835 1.070 ;
        RECT  2.485 0.925 2.605 1.345 ;
        RECT  1.675 1.255 2.485 1.345 ;
        RECT  2.150 0.305 2.260 1.165 ;
        RECT  2.015 0.305 2.150 0.415 ;
        RECT  2.065 1.075 2.150 1.165 ;
        RECT  1.490 0.275 1.705 0.405 ;
        RECT  1.565 0.810 1.675 1.345 ;
        RECT  1.245 0.810 1.565 0.900 ;
        RECT  0.705 0.275 1.490 0.365 ;
        RECT  1.155 0.475 1.245 1.345 ;
        RECT  1.060 0.475 1.155 0.645 ;
        RECT  0.955 1.255 1.155 1.345 ;
        RECT  0.965 0.840 1.065 1.065 ;
        RECT  0.875 0.480 0.965 0.930 ;
        RECT  0.845 1.255 0.955 1.525 ;
        RECT  0.535 0.480 0.875 0.570 ;
        RECT  0.500 0.275 0.705 0.385 ;
        RECT  0.445 0.480 0.535 1.090 ;
        RECT  0.185 0.480 0.445 0.570 ;
        RECT  0.185 1.000 0.445 1.090 ;
        RECT  0.075 0.270 0.185 0.570 ;
        RECT  0.075 1.000 0.185 1.360 ;
    END
END SEDFKCNQD0

MACRO SEDFKCNQD1
    CLASS CORE ;
    FOREIGN SEDFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0203 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.900 2.760 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0580 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.800 3.495 1.120 ;
        RECT  3.350 0.800 3.385 0.890 ;
        RECT  3.045 0.710 3.350 0.890 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.275 7.750 1.490 ;
        RECT  7.620 0.275 7.650 0.675 ;
        RECT  7.620 1.020 7.650 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.190 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.810 1.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.900 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.585 -0.165 7.800 0.165 ;
        RECT  5.585 0.475 5.755 0.585 ;
        RECT  5.485 -0.165 5.585 0.585 ;
        RECT  2.865 -0.165 5.485 0.165 ;
        RECT  2.760 -0.165 2.865 0.600 ;
        RECT  0.000 -0.165 2.760 0.165 ;
        RECT  2.525 0.490 2.760 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.790 1.635 7.800 1.965 ;
        RECT  5.600 1.435 5.790 1.965 ;
        RECT  2.820 1.635 5.600 1.965 ;
        RECT  2.675 1.385 2.820 1.965 ;
        RECT  0.455 1.635 2.675 1.965 ;
        RECT  0.325 1.250 0.455 1.965 ;
        RECT  0.000 1.635 0.325 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.440 0.285 7.530 1.495 ;
        RECT  6.610 0.285 7.440 0.385 ;
        RECT  6.050 1.395 7.440 1.495 ;
        RECT  7.220 0.505 7.330 1.305 ;
        RECT  6.765 0.505 7.220 0.615 ;
        RECT  7.035 1.185 7.220 1.305 ;
        RECT  6.945 0.755 7.020 0.925 ;
        RECT  6.855 0.755 6.945 1.305 ;
        RECT  6.285 1.215 6.855 1.305 ;
        RECT  6.655 0.505 6.765 1.120 ;
        RECT  6.495 0.255 6.610 0.425 ;
        RECT  6.405 0.585 6.515 1.120 ;
        RECT  6.315 0.275 6.405 0.675 ;
        RECT  6.175 0.275 6.315 0.365 ;
        RECT  6.225 0.830 6.285 1.305 ;
        RECT  6.180 0.505 6.225 1.305 ;
        RECT  6.115 0.505 6.180 0.930 ;
        RECT  5.970 0.255 6.175 0.365 ;
        RECT  6.020 1.020 6.090 1.140 ;
        RECT  5.940 1.230 6.050 1.495 ;
        RECT  5.965 0.675 6.020 1.140 ;
        RECT  5.920 0.465 5.965 1.140 ;
        RECT  5.465 1.230 5.940 1.330 ;
        RECT  5.855 0.465 5.920 0.765 ;
        RECT  5.580 0.675 5.855 0.765 ;
        RECT  5.720 0.875 5.830 1.120 ;
        RECT  5.265 1.030 5.720 1.120 ;
        RECT  5.460 0.675 5.580 0.915 ;
        RECT  5.375 1.230 5.465 1.525 ;
        RECT  3.040 1.435 5.375 1.525 ;
        RECT  5.220 1.030 5.265 1.345 ;
        RECT  5.155 0.300 5.220 1.345 ;
        RECT  5.110 0.300 5.155 1.120 ;
        RECT  4.865 1.215 5.050 1.345 ;
        RECT  4.870 0.520 4.985 1.125 ;
        RECT  4.795 0.255 4.965 0.365 ;
        RECT  4.560 0.520 4.870 0.635 ;
        RECT  4.620 1.015 4.870 1.125 ;
        RECT  3.395 1.255 4.865 1.345 ;
        RECT  3.310 0.275 4.795 0.365 ;
        RECT  4.350 0.775 4.645 0.895 ;
        RECT  4.260 0.500 4.350 1.145 ;
        RECT  4.000 0.500 4.260 0.610 ;
        RECT  4.075 1.035 4.260 1.145 ;
        RECT  3.615 0.600 3.725 1.165 ;
        RECT  3.555 0.600 3.615 0.690 ;
        RECT  3.445 0.475 3.555 0.690 ;
        RECT  3.190 1.215 3.395 1.345 ;
        RECT  3.140 0.275 3.310 0.585 ;
        RECT  2.940 0.990 3.240 1.090 ;
        RECT  2.940 1.205 3.040 1.525 ;
        RECT  2.850 0.700 2.940 1.090 ;
        RECT  2.585 1.205 2.940 1.295 ;
        RECT  2.435 0.700 2.850 0.790 ;
        RECT  2.495 1.205 2.585 1.525 ;
        RECT  1.450 1.435 2.495 1.525 ;
        RECT  2.350 0.475 2.435 0.790 ;
        RECT  2.350 1.175 2.405 1.345 ;
        RECT  2.260 0.475 2.350 1.345 ;
        RECT  2.170 0.265 2.290 0.375 ;
        RECT  2.080 0.265 2.170 1.340 ;
        RECT  2.050 0.265 2.080 0.655 ;
        RECT  2.030 1.170 2.080 1.340 ;
        RECT  1.960 0.750 1.990 0.920 ;
        RECT  1.850 0.495 1.960 1.080 ;
        RECT  1.265 0.495 1.850 0.600 ;
        RECT  1.665 0.990 1.850 1.080 ;
        RECT  1.495 0.275 1.705 0.405 ;
        RECT  1.540 0.990 1.665 1.345 ;
        RECT  0.715 0.275 1.495 0.365 ;
        RECT  1.360 1.010 1.450 1.525 ;
        RECT  1.175 0.475 1.265 1.330 ;
        RECT  1.095 0.475 1.175 0.665 ;
        RECT  0.965 1.240 1.175 1.330 ;
        RECT  0.990 0.875 1.085 1.085 ;
        RECT  0.900 0.525 0.990 1.085 ;
        RECT  0.835 1.240 0.965 1.515 ;
        RECT  0.540 0.525 0.900 0.615 ;
        RECT  0.575 0.255 0.715 0.435 ;
        RECT  0.435 0.525 0.540 1.140 ;
        RECT  0.410 0.315 0.435 1.140 ;
        RECT  0.325 0.315 0.410 0.625 ;
        RECT  0.195 1.040 0.410 1.140 ;
        RECT  0.065 1.040 0.195 1.420 ;
    END
END SEDFKCNQD1

MACRO SEDFKCNQD2
    CLASS CORE ;
    FOREIGN SEDFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0203 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.900 2.760 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0580 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.800 3.495 1.120 ;
        RECT  3.350 0.800 3.385 0.890 ;
        RECT  3.045 0.710 3.350 0.890 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.575 7.750 1.120 ;
        RECT  7.645 0.575 7.650 0.675 ;
        RECT  7.645 1.020 7.650 1.120 ;
        RECT  7.535 0.275 7.645 0.675 ;
        RECT  7.535 1.020 7.645 1.425 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.190 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.810 1.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0279 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.900 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.905 -0.165 8.000 0.165 ;
        RECT  7.795 -0.165 7.905 0.485 ;
        RECT  5.525 -0.165 7.795 0.165 ;
        RECT  5.525 0.475 5.695 0.585 ;
        RECT  5.425 -0.165 5.525 0.585 ;
        RECT  2.865 -0.165 5.425 0.165 ;
        RECT  2.760 -0.165 2.865 0.600 ;
        RECT  0.000 -0.165 2.760 0.165 ;
        RECT  2.525 0.490 2.760 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.905 1.635 8.000 1.965 ;
        RECT  7.795 1.220 7.905 1.965 ;
        RECT  5.730 1.635 7.795 1.965 ;
        RECT  5.540 1.435 5.730 1.965 ;
        RECT  2.820 1.635 5.540 1.965 ;
        RECT  2.675 1.385 2.820 1.965 ;
        RECT  0.455 1.635 2.675 1.965 ;
        RECT  0.325 1.250 0.455 1.965 ;
        RECT  0.000 1.635 0.325 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.355 0.285 7.445 1.495 ;
        RECT  6.550 0.285 7.355 0.385 ;
        RECT  5.990 1.395 7.355 1.495 ;
        RECT  7.155 0.755 7.265 0.925 ;
        RECT  7.065 0.505 7.155 1.305 ;
        RECT  6.705 0.505 7.065 0.615 ;
        RECT  6.985 1.115 7.065 1.305 ;
        RECT  6.885 0.755 6.960 0.925 ;
        RECT  6.795 0.755 6.885 1.305 ;
        RECT  6.225 1.215 6.795 1.305 ;
        RECT  6.595 0.505 6.705 1.120 ;
        RECT  6.435 0.255 6.550 0.425 ;
        RECT  6.345 0.585 6.455 1.120 ;
        RECT  6.255 0.275 6.345 0.675 ;
        RECT  6.115 0.275 6.255 0.365 ;
        RECT  6.165 0.830 6.225 1.305 ;
        RECT  6.120 0.505 6.165 1.305 ;
        RECT  6.055 0.505 6.120 0.930 ;
        RECT  5.910 0.255 6.115 0.365 ;
        RECT  5.960 1.020 6.030 1.140 ;
        RECT  5.880 1.230 5.990 1.495 ;
        RECT  5.905 0.675 5.960 1.140 ;
        RECT  5.860 0.465 5.905 1.140 ;
        RECT  5.405 1.230 5.880 1.330 ;
        RECT  5.795 0.465 5.860 0.765 ;
        RECT  5.520 0.675 5.795 0.765 ;
        RECT  5.660 0.875 5.770 1.120 ;
        RECT  5.205 1.030 5.660 1.120 ;
        RECT  5.400 0.675 5.520 0.915 ;
        RECT  5.315 1.230 5.405 1.525 ;
        RECT  3.040 1.435 5.315 1.525 ;
        RECT  5.160 1.030 5.205 1.345 ;
        RECT  5.095 0.300 5.160 1.345 ;
        RECT  5.050 0.300 5.095 1.120 ;
        RECT  4.805 1.215 4.990 1.345 ;
        RECT  4.810 0.520 4.925 1.125 ;
        RECT  4.735 0.255 4.905 0.365 ;
        RECT  4.500 0.520 4.810 0.635 ;
        RECT  4.580 1.015 4.810 1.125 ;
        RECT  3.395 1.255 4.805 1.345 ;
        RECT  3.310 0.275 4.735 0.365 ;
        RECT  4.350 0.775 4.590 0.895 ;
        RECT  4.260 0.500 4.350 1.145 ;
        RECT  4.000 0.500 4.260 0.610 ;
        RECT  4.075 1.035 4.260 1.145 ;
        RECT  3.615 0.600 3.725 1.165 ;
        RECT  3.555 0.600 3.615 0.690 ;
        RECT  3.445 0.475 3.555 0.690 ;
        RECT  3.190 1.215 3.395 1.345 ;
        RECT  3.140 0.275 3.310 0.585 ;
        RECT  2.940 0.990 3.240 1.090 ;
        RECT  2.940 1.205 3.040 1.525 ;
        RECT  2.850 0.700 2.940 1.090 ;
        RECT  2.585 1.205 2.940 1.295 ;
        RECT  2.435 0.700 2.850 0.790 ;
        RECT  2.495 1.205 2.585 1.525 ;
        RECT  1.450 1.435 2.495 1.525 ;
        RECT  2.350 0.475 2.435 0.790 ;
        RECT  2.350 1.175 2.405 1.345 ;
        RECT  2.260 0.475 2.350 1.345 ;
        RECT  2.170 0.265 2.290 0.375 ;
        RECT  2.080 0.265 2.170 1.340 ;
        RECT  2.050 0.265 2.080 0.655 ;
        RECT  2.030 1.170 2.080 1.340 ;
        RECT  1.960 0.750 1.990 0.920 ;
        RECT  1.850 0.495 1.960 1.080 ;
        RECT  1.265 0.495 1.850 0.600 ;
        RECT  1.665 0.990 1.850 1.080 ;
        RECT  1.495 0.275 1.705 0.405 ;
        RECT  1.540 0.990 1.665 1.345 ;
        RECT  0.715 0.275 1.495 0.365 ;
        RECT  1.360 1.010 1.450 1.525 ;
        RECT  1.175 0.475 1.265 1.330 ;
        RECT  1.095 0.475 1.175 0.665 ;
        RECT  0.965 1.240 1.175 1.330 ;
        RECT  0.990 0.875 1.085 1.085 ;
        RECT  0.900 0.525 0.990 1.085 ;
        RECT  0.835 1.240 0.965 1.515 ;
        RECT  0.540 0.525 0.900 0.615 ;
        RECT  0.575 0.255 0.715 0.435 ;
        RECT  0.435 0.525 0.540 1.140 ;
        RECT  0.410 0.315 0.435 1.140 ;
        RECT  0.325 0.315 0.410 0.625 ;
        RECT  0.195 1.040 0.410 1.140 ;
        RECT  0.065 1.040 0.195 1.420 ;
    END
END SEDFKCNQD2

MACRO SEDFKCNQD4
    CLASS CORE ;
    FOREIGN SEDFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0203 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.900 2.760 1.090 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0580 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.800 3.495 1.120 ;
        RECT  3.350 0.800 3.385 0.890 ;
        RECT  3.045 0.710 3.350 0.890 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 0.510 8.105 0.690 ;
        RECT  7.850 1.110 8.105 1.290 ;
        RECT  7.550 0.510 7.850 1.290 ;
        RECT  7.435 0.510 7.550 0.690 ;
        RECT  7.435 1.110 7.550 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.190 0.920 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0431 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.810 1.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0551 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.710 4.150 0.890 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0446 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.750 0.900 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.505 -0.165 8.400 0.165 ;
        RECT  5.505 0.475 5.675 0.585 ;
        RECT  5.405 -0.165 5.505 0.585 ;
        RECT  2.865 -0.165 5.405 0.165 ;
        RECT  2.760 -0.165 2.865 0.600 ;
        RECT  0.000 -0.165 2.760 0.165 ;
        RECT  2.525 0.490 2.760 0.600 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.710 1.635 8.400 1.965 ;
        RECT  5.520 1.435 5.710 1.965 ;
        RECT  2.820 1.635 5.520 1.965 ;
        RECT  2.675 1.385 2.820 1.965 ;
        RECT  0.455 1.635 2.675 1.965 ;
        RECT  0.325 1.250 0.455 1.965 ;
        RECT  0.000 1.635 0.325 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.950 0.510 8.105 0.690 ;
        RECT  7.950 1.110 8.105 1.290 ;
        RECT  7.435 0.510 7.450 0.690 ;
        RECT  7.435 1.110 7.450 1.290 ;
        RECT  8.195 0.285 8.285 1.495 ;
        RECT  6.530 0.285 8.195 0.385 ;
        RECT  5.970 1.395 8.195 1.495 ;
        RECT  7.300 0.785 7.440 0.895 ;
        RECT  7.210 0.505 7.300 1.305 ;
        RECT  6.685 0.505 7.210 0.615 ;
        RECT  6.965 1.115 7.210 1.305 ;
        RECT  6.865 0.785 7.080 0.895 ;
        RECT  6.775 0.785 6.865 1.305 ;
        RECT  6.205 1.215 6.775 1.305 ;
        RECT  6.575 0.505 6.685 1.120 ;
        RECT  6.415 0.255 6.530 0.425 ;
        RECT  6.325 0.585 6.435 1.120 ;
        RECT  6.235 0.275 6.325 0.675 ;
        RECT  6.095 0.275 6.235 0.365 ;
        RECT  6.145 0.830 6.205 1.305 ;
        RECT  6.100 0.505 6.145 1.305 ;
        RECT  6.035 0.505 6.100 0.930 ;
        RECT  5.890 0.255 6.095 0.365 ;
        RECT  5.940 1.020 6.010 1.140 ;
        RECT  5.860 1.230 5.970 1.495 ;
        RECT  5.885 0.675 5.940 1.140 ;
        RECT  5.840 0.465 5.885 1.140 ;
        RECT  5.385 1.230 5.860 1.330 ;
        RECT  5.775 0.465 5.840 0.765 ;
        RECT  5.500 0.675 5.775 0.765 ;
        RECT  5.640 0.875 5.750 1.120 ;
        RECT  5.185 1.030 5.640 1.120 ;
        RECT  5.380 0.675 5.500 0.915 ;
        RECT  5.295 1.230 5.385 1.525 ;
        RECT  3.040 1.435 5.295 1.525 ;
        RECT  5.140 1.030 5.185 1.345 ;
        RECT  5.075 0.300 5.140 1.345 ;
        RECT  5.030 0.300 5.075 1.120 ;
        RECT  4.785 1.215 4.970 1.345 ;
        RECT  4.790 0.520 4.905 1.125 ;
        RECT  4.715 0.255 4.885 0.365 ;
        RECT  4.500 0.520 4.790 0.635 ;
        RECT  4.540 1.015 4.790 1.125 ;
        RECT  3.395 1.255 4.785 1.345 ;
        RECT  3.310 0.275 4.715 0.365 ;
        RECT  4.350 0.775 4.590 0.895 ;
        RECT  4.260 0.500 4.350 1.145 ;
        RECT  4.000 0.500 4.260 0.610 ;
        RECT  4.075 1.035 4.260 1.145 ;
        RECT  3.615 0.600 3.725 1.165 ;
        RECT  3.555 0.600 3.615 0.690 ;
        RECT  3.445 0.475 3.555 0.690 ;
        RECT  3.190 1.215 3.395 1.345 ;
        RECT  3.140 0.275 3.310 0.585 ;
        RECT  2.940 0.990 3.240 1.090 ;
        RECT  2.940 1.205 3.040 1.525 ;
        RECT  2.850 0.700 2.940 1.090 ;
        RECT  2.585 1.205 2.940 1.295 ;
        RECT  2.435 0.700 2.850 0.790 ;
        RECT  2.495 1.205 2.585 1.525 ;
        RECT  1.450 1.435 2.495 1.525 ;
        RECT  2.350 0.475 2.435 0.790 ;
        RECT  2.350 1.175 2.405 1.345 ;
        RECT  2.260 0.475 2.350 1.345 ;
        RECT  2.170 0.265 2.290 0.375 ;
        RECT  2.080 0.265 2.170 1.340 ;
        RECT  2.050 0.265 2.080 0.655 ;
        RECT  2.030 1.170 2.080 1.340 ;
        RECT  1.960 0.750 1.990 0.920 ;
        RECT  1.850 0.495 1.960 1.080 ;
        RECT  1.265 0.495 1.850 0.600 ;
        RECT  1.665 0.990 1.850 1.080 ;
        RECT  1.495 0.275 1.705 0.405 ;
        RECT  1.540 0.990 1.665 1.345 ;
        RECT  0.715 0.275 1.495 0.365 ;
        RECT  1.360 1.010 1.450 1.525 ;
        RECT  1.175 0.475 1.265 1.330 ;
        RECT  1.095 0.475 1.175 0.665 ;
        RECT  0.965 1.240 1.175 1.330 ;
        RECT  0.990 0.875 1.085 1.085 ;
        RECT  0.900 0.525 0.990 1.085 ;
        RECT  0.835 1.240 0.965 1.515 ;
        RECT  0.540 0.525 0.900 0.615 ;
        RECT  0.575 0.255 0.715 0.435 ;
        RECT  0.435 0.525 0.540 1.140 ;
        RECT  0.410 0.315 0.435 1.140 ;
        RECT  0.325 0.315 0.410 0.625 ;
        RECT  0.195 1.040 0.410 1.140 ;
        RECT  0.065 1.040 0.195 1.420 ;
    END
END SEDFKCNQD4

MACRO SEDFQD0
    CLASS CORE ;
    FOREIGN SEDFQD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0710 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.340 6.350 1.545 ;
        RECT  6.135 0.340 6.250 0.450 ;
        RECT  6.165 1.335 6.250 1.545 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0495 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 -0.165 6.600 0.165 ;
        RECT  5.620 -0.165 5.730 0.450 ;
        RECT  2.110 -0.165 5.620 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 6.600 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.070 0.560 6.160 1.120 ;
        RECT  6.015 0.560 6.070 0.670 ;
        RECT  5.960 1.010 6.070 1.525 ;
        RECT  5.905 0.425 6.015 0.670 ;
        RECT  5.855 0.780 5.960 0.890 ;
        RECT  5.000 1.435 5.960 1.525 ;
        RECT  5.665 0.560 5.905 0.670 ;
        RECT  5.765 0.780 5.855 1.345 ;
        RECT  5.205 1.255 5.765 1.345 ;
        RECT  5.555 0.560 5.665 0.920 ;
        RECT  5.465 1.060 5.525 1.165 ;
        RECT  5.375 0.275 5.465 1.165 ;
        RECT  5.160 0.275 5.375 0.365 ;
        RECT  5.350 1.060 5.375 1.165 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.990 0.255 5.160 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.990 0.365 ;
        RECT  4.885 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.795 0.735 4.845 0.905 ;
        RECT  4.705 0.475 4.795 0.905 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.750 3.655 0.920 ;
        RECT  3.440 0.515 3.530 1.165 ;
        RECT  3.135 0.515 3.440 0.620 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.305 0.360 1.090 ;
        RECT  0.045 0.305 0.270 0.415 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQD0

MACRO SEDFQD1
    CLASS CORE ;
    FOREIGN SEDFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1350 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.340 6.350 1.490 ;
        RECT  6.135 0.340 6.250 0.450 ;
        RECT  6.165 1.280 6.250 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.735 -0.165 6.600 0.165 ;
        RECT  5.625 -0.165 5.735 0.450 ;
        RECT  2.110 -0.165 5.625 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 6.600 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.070 0.560 6.160 1.120 ;
        RECT  6.020 0.560 6.070 0.670 ;
        RECT  5.960 1.010 6.070 1.525 ;
        RECT  5.910 0.425 6.020 0.670 ;
        RECT  5.855 0.780 5.960 0.890 ;
        RECT  5.000 1.435 5.960 1.525 ;
        RECT  5.665 0.560 5.910 0.670 ;
        RECT  5.765 0.780 5.855 1.345 ;
        RECT  5.205 1.255 5.765 1.345 ;
        RECT  5.555 0.560 5.665 0.920 ;
        RECT  5.465 1.060 5.525 1.165 ;
        RECT  5.375 0.275 5.465 1.165 ;
        RECT  5.160 0.275 5.375 0.365 ;
        RECT  5.350 1.060 5.375 1.165 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.990 0.255 5.160 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.990 0.365 ;
        RECT  4.885 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.795 0.735 4.845 0.905 ;
        RECT  4.705 0.475 4.795 0.905 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.740 3.655 0.910 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQD1

MACRO SEDFQD2
    CLASS CORE ;
    FOREIGN SEDFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.565 6.750 1.180 ;
        RECT  6.615 0.565 6.650 0.665 ;
        RECT  6.615 1.080 6.650 1.180 ;
        RECT  6.505 0.295 6.615 0.665 ;
        RECT  6.505 1.080 6.615 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.875 -0.165 7.000 0.165 ;
        RECT  6.765 -0.165 6.875 0.465 ;
        RECT  6.355 -0.165 6.765 0.165 ;
        RECT  6.245 -0.165 6.355 0.465 ;
        RECT  5.735 -0.165 6.245 0.165 ;
        RECT  5.625 -0.165 5.735 0.450 ;
        RECT  2.110 -0.165 5.625 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.875 1.635 7.000 1.965 ;
        RECT  6.765 1.280 6.875 1.965 ;
        RECT  6.355 1.635 6.765 1.965 ;
        RECT  6.250 1.280 6.355 1.965 ;
        RECT  4.740 1.635 6.250 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.305 0.560 6.395 1.120 ;
        RECT  6.020 0.560 6.305 0.670 ;
        RECT  6.070 1.010 6.305 1.120 ;
        RECT  5.855 0.780 6.165 0.890 ;
        RECT  5.960 1.010 6.070 1.525 ;
        RECT  5.910 0.425 6.020 0.670 ;
        RECT  5.000 1.435 5.960 1.525 ;
        RECT  5.665 0.560 5.910 0.670 ;
        RECT  5.765 0.780 5.855 1.345 ;
        RECT  5.205 1.255 5.765 1.345 ;
        RECT  5.555 0.560 5.665 0.920 ;
        RECT  5.465 1.060 5.525 1.165 ;
        RECT  5.375 0.275 5.465 1.165 ;
        RECT  5.160 0.275 5.375 0.365 ;
        RECT  5.350 1.060 5.375 1.165 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.990 0.255 5.160 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.990 0.365 ;
        RECT  4.885 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.795 0.735 4.845 0.905 ;
        RECT  4.705 0.475 4.795 0.905 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.740 3.655 0.910 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQD2

MACRO SEDFQD4
    CLASS CORE ;
    FOREIGN SEDFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.325 7.695 0.635 ;
        RECT  7.450 1.100 7.695 1.410 ;
        RECT  7.150 0.325 7.450 1.410 ;
        RECT  7.015 0.325 7.150 0.635 ;
        RECT  7.015 1.100 7.150 1.410 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.895 -0.165 8.000 0.165 ;
        RECT  6.785 -0.165 6.895 0.450 ;
        RECT  6.335 -0.165 6.785 0.165 ;
        RECT  6.225 -0.165 6.335 0.450 ;
        RECT  2.110 -0.165 6.225 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.895 1.635 8.000 1.965 ;
        RECT  6.785 1.350 6.895 1.965 ;
        RECT  5.330 1.635 6.785 1.965 ;
        RECT  5.160 1.445 5.330 1.965 ;
        RECT  4.760 1.635 5.160 1.965 ;
        RECT  4.590 1.445 4.760 1.965 ;
        RECT  0.525 1.635 4.590 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.550 0.325 7.695 0.635 ;
        RECT  7.550 1.100 7.695 1.410 ;
        RECT  7.015 0.325 7.050 0.635 ;
        RECT  7.015 1.100 7.050 1.410 ;
        RECT  6.835 0.560 6.925 1.120 ;
        RECT  6.620 0.560 6.835 0.670 ;
        RECT  6.670 1.010 6.835 1.120 ;
        RECT  6.455 0.780 6.745 0.890 ;
        RECT  6.560 1.010 6.670 1.525 ;
        RECT  6.510 0.425 6.620 0.670 ;
        RECT  5.600 1.435 6.560 1.525 ;
        RECT  6.265 0.560 6.510 0.670 ;
        RECT  6.365 0.780 6.455 1.345 ;
        RECT  5.805 1.255 6.365 1.345 ;
        RECT  6.155 0.560 6.265 0.920 ;
        RECT  6.065 1.060 6.125 1.165 ;
        RECT  5.975 0.275 6.065 1.165 ;
        RECT  5.760 0.275 5.975 0.365 ;
        RECT  5.950 1.060 5.975 1.165 ;
        RECT  5.805 0.465 5.885 0.575 ;
        RECT  5.715 0.465 5.805 1.345 ;
        RECT  5.590 0.255 5.760 0.365 ;
        RECT  5.450 0.485 5.625 1.155 ;
        RECT  5.510 1.265 5.600 1.525 ;
        RECT  4.435 0.275 5.590 0.365 ;
        RECT  4.335 1.265 5.510 1.355 ;
        RECT  4.880 0.485 5.450 0.595 ;
        RECT  4.610 1.045 5.450 1.155 ;
        RECT  4.790 0.765 5.010 0.875 ;
        RECT  4.700 0.475 4.790 0.875 ;
        RECT  4.365 0.475 4.700 0.565 ;
        RECT  4.510 0.710 4.610 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.245 1.265 4.335 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.125 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.245 1.525 ;
        RECT  3.845 0.725 4.110 0.835 ;
        RECT  3.835 1.235 4.040 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  2.495 1.255 3.835 1.345 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.750 3.655 0.920 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQD4

MACRO SEDFQND0
    CLASS CORE ;
    FOREIGN SEDFQND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0710 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.340 6.350 1.545 ;
        RECT  6.135 0.340 6.250 0.450 ;
        RECT  6.165 1.335 6.250 1.545 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0495 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 -0.165 6.600 0.165 ;
        RECT  5.620 -0.165 5.730 0.450 ;
        RECT  2.110 -0.165 5.620 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 6.600 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.070 0.560 6.160 1.120 ;
        RECT  6.060 0.560 6.070 1.525 ;
        RECT  6.015 0.560 6.060 0.670 ;
        RECT  5.960 1.010 6.060 1.525 ;
        RECT  5.905 0.425 6.015 0.670 ;
        RECT  5.000 1.435 5.960 1.525 ;
        RECT  5.855 0.780 5.955 0.890 ;
        RECT  5.665 0.560 5.905 0.670 ;
        RECT  5.765 0.780 5.855 1.345 ;
        RECT  5.205 1.255 5.765 1.345 ;
        RECT  5.555 0.560 5.665 0.920 ;
        RECT  5.465 1.060 5.525 1.165 ;
        RECT  5.375 0.275 5.465 1.165 ;
        RECT  5.160 0.275 5.375 0.365 ;
        RECT  5.350 1.060 5.375 1.165 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.990 0.255 5.160 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.990 0.365 ;
        RECT  4.885 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.795 0.735 4.845 0.905 ;
        RECT  4.705 0.475 4.795 0.905 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.750 3.655 0.920 ;
        RECT  3.440 0.515 3.530 1.165 ;
        RECT  3.135 0.515 3.440 0.620 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.305 0.360 1.090 ;
        RECT  0.045 0.305 0.270 0.415 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQND0

MACRO SEDFQND1
    CLASS CORE ;
    FOREIGN SEDFQND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1350 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 0.340 6.350 1.490 ;
        RECT  6.135 0.340 6.250 0.450 ;
        RECT  6.165 1.280 6.250 1.490 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.735 -0.165 6.600 0.165 ;
        RECT  5.625 -0.165 5.735 0.450 ;
        RECT  2.110 -0.165 5.625 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 6.600 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.070 0.560 6.160 1.120 ;
        RECT  6.060 0.560 6.070 1.525 ;
        RECT  6.020 0.560 6.060 0.670 ;
        RECT  5.960 1.010 6.060 1.525 ;
        RECT  5.910 0.425 6.020 0.670 ;
        RECT  5.855 0.780 5.960 0.890 ;
        RECT  5.000 1.435 5.960 1.525 ;
        RECT  5.665 0.560 5.910 0.670 ;
        RECT  5.765 0.780 5.855 1.345 ;
        RECT  5.205 1.255 5.765 1.345 ;
        RECT  5.555 0.560 5.665 0.920 ;
        RECT  5.465 1.060 5.525 1.165 ;
        RECT  5.375 0.275 5.465 1.165 ;
        RECT  5.160 0.275 5.375 0.365 ;
        RECT  5.350 1.060 5.375 1.165 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.990 0.255 5.160 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.990 0.365 ;
        RECT  4.885 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.795 0.735 4.845 0.905 ;
        RECT  4.705 0.475 4.795 0.905 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.740 3.655 0.910 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQND1

MACRO SEDFQND2
    CLASS CORE ;
    FOREIGN SEDFQND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.650 0.565 6.750 1.180 ;
        RECT  6.615 0.565 6.650 0.665 ;
        RECT  6.615 1.080 6.650 1.180 ;
        RECT  6.505 0.295 6.615 0.665 ;
        RECT  6.505 1.080 6.615 1.490 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0282 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.875 -0.165 7.000 0.165 ;
        RECT  6.765 -0.165 6.875 0.465 ;
        RECT  6.355 -0.165 6.765 0.165 ;
        RECT  6.245 -0.165 6.355 0.465 ;
        RECT  5.735 -0.165 6.245 0.165 ;
        RECT  5.625 -0.165 5.735 0.450 ;
        RECT  2.110 -0.165 5.625 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.875 1.635 7.000 1.965 ;
        RECT  6.765 1.280 6.875 1.965 ;
        RECT  6.355 1.635 6.765 1.965 ;
        RECT  6.250 1.280 6.355 1.965 ;
        RECT  4.740 1.635 6.250 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.285 0.560 6.395 1.120 ;
        RECT  6.020 0.560 6.285 0.670 ;
        RECT  6.070 1.010 6.285 1.120 ;
        RECT  5.960 1.010 6.070 1.525 ;
        RECT  5.910 0.425 6.020 0.670 ;
        RECT  5.855 0.780 5.965 0.890 ;
        RECT  5.000 1.435 5.960 1.525 ;
        RECT  5.665 0.560 5.910 0.670 ;
        RECT  5.765 0.780 5.855 1.345 ;
        RECT  5.205 1.255 5.765 1.345 ;
        RECT  5.555 0.560 5.665 0.920 ;
        RECT  5.465 1.060 5.525 1.165 ;
        RECT  5.375 0.275 5.465 1.165 ;
        RECT  5.160 0.275 5.375 0.365 ;
        RECT  5.350 1.060 5.375 1.165 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.990 0.255 5.160 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.990 0.365 ;
        RECT  4.885 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.795 0.735 4.845 0.905 ;
        RECT  4.705 0.475 4.795 0.905 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.740 3.655 0.910 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQND2

MACRO SEDFQND4
    CLASS CORE ;
    FOREIGN SEDFQND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0190 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.510 1.550 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.685 2.950 1.090 ;
        RECT  2.555 0.685 2.840 0.785 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.325 7.105 0.635 ;
        RECT  6.850 1.100 7.105 1.410 ;
        RECT  6.550 0.325 6.850 1.410 ;
        RECT  6.435 0.325 6.550 0.635 ;
        RECT  6.435 1.100 6.550 1.410 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0554 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.510 0.180 0.890 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0277 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.760 0.700 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.710 3.350 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.295 -0.165 7.400 0.165 ;
        RECT  6.185 -0.165 6.295 0.450 ;
        RECT  5.735 -0.165 6.185 0.165 ;
        RECT  5.625 -0.165 5.735 0.450 ;
        RECT  2.110 -0.165 5.625 0.165 ;
        RECT  2.000 -0.165 2.110 0.395 ;
        RECT  0.000 -0.165 2.000 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 1.635 7.400 1.965 ;
        RECT  4.570 1.445 4.740 1.965 ;
        RECT  0.525 1.635 4.570 1.965 ;
        RECT  0.435 1.180 0.525 1.965 ;
        RECT  0.300 1.180 0.435 1.290 ;
        RECT  0.000 1.635 0.435 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.950 0.325 7.105 0.635 ;
        RECT  6.950 1.100 7.105 1.410 ;
        RECT  6.435 0.325 6.450 0.635 ;
        RECT  6.435 1.100 6.450 1.410 ;
        RECT  6.210 0.750 6.415 0.920 ;
        RECT  6.110 0.560 6.210 1.120 ;
        RECT  6.020 0.560 6.110 0.670 ;
        RECT  6.070 1.010 6.110 1.120 ;
        RECT  5.960 1.010 6.070 1.525 ;
        RECT  5.910 0.295 6.020 0.670 ;
        RECT  5.000 1.435 5.960 1.525 ;
        RECT  5.855 0.780 5.955 0.890 ;
        RECT  5.665 0.560 5.910 0.670 ;
        RECT  5.765 0.780 5.855 1.345 ;
        RECT  5.205 1.255 5.765 1.345 ;
        RECT  5.555 0.560 5.665 0.920 ;
        RECT  5.465 1.060 5.525 1.165 ;
        RECT  5.375 0.275 5.465 1.165 ;
        RECT  5.160 0.275 5.375 0.365 ;
        RECT  5.350 1.060 5.375 1.165 ;
        RECT  5.205 0.465 5.285 0.575 ;
        RECT  5.115 0.465 5.205 1.345 ;
        RECT  4.990 0.255 5.160 0.365 ;
        RECT  4.935 0.455 5.025 1.155 ;
        RECT  4.910 1.265 5.000 1.525 ;
        RECT  4.435 0.275 4.990 0.365 ;
        RECT  4.885 0.455 4.935 0.645 ;
        RECT  4.615 1.045 4.935 1.155 ;
        RECT  4.340 1.265 4.910 1.355 ;
        RECT  4.795 0.735 4.845 0.905 ;
        RECT  4.705 0.475 4.795 0.905 ;
        RECT  4.365 0.475 4.705 0.565 ;
        RECT  4.515 0.710 4.615 1.155 ;
        RECT  4.265 0.255 4.435 0.365 ;
        RECT  4.275 0.475 4.365 1.175 ;
        RECT  4.250 1.265 4.340 1.525 ;
        RECT  4.145 0.475 4.275 0.575 ;
        RECT  4.130 1.065 4.275 1.175 ;
        RECT  1.100 1.435 4.250 1.525 ;
        RECT  3.845 0.725 4.115 0.835 ;
        RECT  3.840 1.235 4.045 1.345 ;
        RECT  3.835 0.255 4.005 0.365 ;
        RECT  3.750 0.515 3.845 1.135 ;
        RECT  2.495 1.255 3.840 1.345 ;
        RECT  2.640 0.275 3.835 0.365 ;
        RECT  3.635 0.515 3.750 0.625 ;
        RECT  3.640 1.025 3.750 1.135 ;
        RECT  3.530 0.750 3.655 0.920 ;
        RECT  3.440 0.480 3.530 1.165 ;
        RECT  3.135 0.480 3.440 0.590 ;
        RECT  3.150 1.055 3.440 1.165 ;
        RECT  2.845 0.495 3.015 0.595 ;
        RECT  1.910 0.495 2.845 0.585 ;
        RECT  2.625 0.875 2.730 1.150 ;
        RECT  2.470 0.275 2.640 0.405 ;
        RECT  2.385 0.875 2.625 0.965 ;
        RECT  2.385 1.055 2.515 1.165 ;
        RECT  2.295 0.685 2.385 0.965 ;
        RECT  2.295 1.055 2.385 1.345 ;
        RECT  1.955 0.685 2.295 0.795 ;
        RECT  1.160 1.255 2.295 1.345 ;
        RECT  1.860 0.685 1.955 1.165 ;
        RECT  1.820 0.305 1.910 0.585 ;
        RECT  1.730 0.685 1.860 0.795 ;
        RECT  1.765 1.050 1.860 1.165 ;
        RECT  1.340 0.305 1.820 0.415 ;
        RECT  1.640 0.525 1.730 0.795 ;
        RECT  1.340 1.055 1.675 1.165 ;
        RECT  1.250 0.305 1.340 1.165 ;
        RECT  1.070 0.310 1.160 1.345 ;
        RECT  0.715 0.310 1.070 0.420 ;
        RECT  0.745 1.140 1.070 1.250 ;
        RECT  0.870 0.515 0.980 0.965 ;
        RECT  0.360 0.855 0.870 0.965 ;
        RECT  0.270 0.310 0.360 1.090 ;
        RECT  0.045 0.310 0.270 0.420 ;
        RECT  0.185 1.000 0.270 1.090 ;
        RECT  0.075 1.000 0.185 1.300 ;
    END
END SEDFQND4

MACRO SEDFQNXD0
    CLASS CORE ;
    FOREIGN SEDFQNXD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.550 0.545 6.845 0.655 ;
        RECT  6.550 1.030 6.845 1.140 ;
        RECT  6.450 0.545 6.550 1.140 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0724 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 7.400 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.460 1.635 7.400 1.965 ;
        RECT  5.290 1.445 5.460 1.965 ;
        RECT  4.930 1.635 5.290 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.265 0.275 7.355 1.525 ;
        RECT  6.315 0.275 7.265 0.365 ;
        RECT  6.310 1.435 7.265 1.525 ;
        RECT  6.645 1.245 7.155 1.345 ;
        RECT  6.965 0.515 7.075 1.155 ;
        RECT  6.650 0.780 6.965 0.890 ;
        RECT  6.555 1.230 6.645 1.345 ;
        RECT  5.925 1.230 6.555 1.320 ;
        RECT  6.215 0.275 6.315 0.645 ;
        RECT  6.140 1.410 6.310 1.525 ;
        RECT  6.125 1.000 6.240 1.110 ;
        RECT  5.720 1.435 6.140 1.525 ;
        RECT  6.035 0.275 6.125 1.110 ;
        RECT  5.875 0.275 6.035 0.365 ;
        RECT  5.925 0.475 5.945 0.645 ;
        RECT  5.835 0.475 5.925 1.320 ;
        RECT  5.705 0.255 5.875 0.365 ;
        RECT  5.655 0.455 5.745 1.155 ;
        RECT  5.630 1.265 5.720 1.525 ;
        RECT  5.140 0.275 5.705 0.365 ;
        RECT  5.595 0.455 5.655 0.645 ;
        RECT  5.320 1.045 5.655 1.155 ;
        RECT  4.650 1.265 5.630 1.355 ;
        RECT  5.500 0.735 5.565 0.905 ;
        RECT  5.410 0.475 5.500 0.905 ;
        RECT  5.120 0.475 5.410 0.565 ;
        RECT  5.220 0.735 5.320 1.155 ;
        RECT  4.970 0.255 5.140 0.365 ;
        RECT  5.030 0.475 5.120 1.175 ;
        RECT  4.855 0.475 5.030 0.575 ;
        RECT  4.855 1.065 5.030 1.175 ;
        RECT  4.585 0.275 4.970 0.365 ;
        RECT  4.765 0.700 4.940 0.810 ;
        RECT  4.675 0.700 4.765 1.175 ;
        RECT  4.470 1.085 4.675 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.475 0.275 4.585 0.995 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.305 0.275 4.475 0.365 ;
        RECT  4.290 0.905 4.475 0.995 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.205 0.275 4.305 0.490 ;
        RECT  4.180 0.905 4.290 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.660 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.190 0.275 3.440 0.415 ;
        RECT  3.305 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.305 1.345 ;
        RECT  3.195 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.195 0.610 ;
        RECT  2.610 1.045 3.195 1.135 ;
        RECT  1.700 0.275 3.190 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQNXD0

MACRO SEDFQNXD1
    CLASS CORE ;
    FOREIGN SEDFQNXD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.550 0.505 6.860 0.615 ;
        RECT  6.550 1.030 6.860 1.140 ;
        RECT  6.450 0.505 6.550 1.140 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 7.400 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.475 1.635 7.400 1.965 ;
        RECT  5.305 1.445 5.475 1.965 ;
        RECT  4.930 1.635 5.305 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.265 0.275 7.355 1.525 ;
        RECT  6.330 0.275 7.265 0.365 ;
        RECT  6.325 1.435 7.265 1.525 ;
        RECT  6.660 1.245 7.155 1.345 ;
        RECT  6.965 0.515 7.075 1.155 ;
        RECT  6.660 0.780 6.965 0.890 ;
        RECT  6.570 1.230 6.660 1.345 ;
        RECT  5.940 1.230 6.570 1.320 ;
        RECT  6.230 0.275 6.330 0.645 ;
        RECT  6.155 1.410 6.325 1.525 ;
        RECT  6.140 1.000 6.255 1.110 ;
        RECT  5.735 1.435 6.155 1.525 ;
        RECT  6.050 0.275 6.140 1.110 ;
        RECT  5.890 0.275 6.050 0.365 ;
        RECT  5.940 0.475 5.960 0.645 ;
        RECT  5.850 0.475 5.940 1.320 ;
        RECT  5.720 0.255 5.890 0.365 ;
        RECT  5.670 0.455 5.760 1.155 ;
        RECT  5.645 1.265 5.735 1.525 ;
        RECT  5.155 0.275 5.720 0.365 ;
        RECT  5.610 0.455 5.670 0.645 ;
        RECT  5.335 1.045 5.670 1.155 ;
        RECT  4.650 1.265 5.645 1.355 ;
        RECT  5.515 0.735 5.580 0.905 ;
        RECT  5.425 0.475 5.515 0.905 ;
        RECT  5.135 0.475 5.425 0.565 ;
        RECT  5.235 0.735 5.335 1.155 ;
        RECT  4.985 0.255 5.155 0.365 ;
        RECT  5.045 0.475 5.135 1.175 ;
        RECT  4.870 0.475 5.045 0.575 ;
        RECT  4.870 1.065 5.045 1.175 ;
        RECT  4.600 0.275 4.985 0.365 ;
        RECT  4.780 0.700 4.940 0.810 ;
        RECT  4.690 0.700 4.780 1.175 ;
        RECT  4.470 1.085 4.690 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.490 0.275 4.600 0.995 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.220 0.275 4.490 0.470 ;
        RECT  4.290 0.905 4.490 0.995 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.180 0.905 4.290 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.675 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.205 0.275 3.440 0.415 ;
        RECT  3.320 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.320 1.345 ;
        RECT  3.210 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.210 0.610 ;
        RECT  2.610 1.045 3.210 1.135 ;
        RECT  1.700 0.275 3.205 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQNXD1

MACRO SEDFQNXD2
    CLASS CORE ;
    FOREIGN SEDFQNXD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.150 0.475 7.275 0.645 ;
        RECT  7.150 1.130 7.275 1.300 ;
        RECT  7.050 0.475 7.150 1.300 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 7.600 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.445 1.635 7.600 1.965 ;
        RECT  5.275 1.445 5.445 1.965 ;
        RECT  4.930 1.635 5.275 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.385 0.275 7.475 1.525 ;
        RECT  6.300 0.275 7.385 0.365 ;
        RECT  6.295 1.435 7.385 1.525 ;
        RECT  6.850 0.505 6.960 1.270 ;
        RECT  6.500 0.505 6.850 0.615 ;
        RECT  6.655 1.160 6.850 1.270 ;
        RECT  6.590 0.750 6.700 1.070 ;
        RECT  6.530 0.980 6.590 1.070 ;
        RECT  6.440 0.980 6.530 1.305 ;
        RECT  6.410 0.505 6.500 0.890 ;
        RECT  5.910 1.205 6.440 1.305 ;
        RECT  6.315 0.780 6.410 0.890 ;
        RECT  6.200 0.275 6.300 0.645 ;
        RECT  6.125 1.395 6.295 1.525 ;
        RECT  6.110 1.005 6.245 1.115 ;
        RECT  5.705 1.435 6.125 1.525 ;
        RECT  6.020 0.275 6.110 1.115 ;
        RECT  5.860 0.275 6.020 0.365 ;
        RECT  5.910 0.475 5.930 0.645 ;
        RECT  5.820 0.475 5.910 1.305 ;
        RECT  5.690 0.255 5.860 0.365 ;
        RECT  5.640 0.455 5.730 1.155 ;
        RECT  5.615 1.265 5.705 1.525 ;
        RECT  5.130 0.275 5.690 0.365 ;
        RECT  5.580 0.455 5.640 0.645 ;
        RECT  5.310 1.045 5.640 1.155 ;
        RECT  4.650 1.265 5.615 1.355 ;
        RECT  5.490 0.735 5.550 0.905 ;
        RECT  5.400 0.475 5.490 0.905 ;
        RECT  5.105 0.475 5.400 0.565 ;
        RECT  5.210 0.735 5.310 1.155 ;
        RECT  4.960 0.255 5.130 0.365 ;
        RECT  5.015 0.475 5.105 1.175 ;
        RECT  4.845 0.475 5.015 0.575 ;
        RECT  4.845 1.065 5.015 1.175 ;
        RECT  4.575 0.275 4.960 0.365 ;
        RECT  4.755 0.700 4.910 0.810 ;
        RECT  4.665 0.700 4.755 1.175 ;
        RECT  4.470 1.085 4.665 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.465 0.275 4.575 0.995 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  4.300 0.275 4.465 0.365 ;
        RECT  4.290 0.905 4.465 0.995 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.190 0.275 4.300 0.490 ;
        RECT  4.180 0.905 4.290 1.165 ;
        RECT  4.080 0.625 4.185 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.650 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.175 0.275 3.440 0.415 ;
        RECT  3.290 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.290 1.345 ;
        RECT  3.180 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.180 0.610 ;
        RECT  2.610 1.045 3.180 1.135 ;
        RECT  1.700 0.275 3.175 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQNXD2

MACRO SEDFQNXD4
    CLASS CORE ;
    FOREIGN SEDFQNXD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.510 7.905 0.690 ;
        RECT  7.650 1.115 7.905 1.285 ;
        RECT  7.350 0.510 7.650 1.285 ;
        RECT  7.235 0.510 7.350 0.690 ;
        RECT  7.235 1.115 7.350 1.285 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0493 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.580 -0.165 8.200 0.165 ;
        RECT  4.470 -0.165 4.580 0.490 ;
        RECT  1.310 -0.165 4.470 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.635 8.200 1.965 ;
        RECT  5.350 1.445 5.520 1.965 ;
        RECT  4.920 1.635 5.350 1.965 ;
        RECT  4.750 1.445 4.920 1.965 ;
        RECT  2.990 1.635 4.750 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.750 0.510 7.905 0.690 ;
        RECT  7.750 1.115 7.905 1.285 ;
        RECT  7.235 0.510 7.250 0.690 ;
        RECT  7.235 1.115 7.250 1.285 ;
        RECT  8.000 0.275 8.090 1.525 ;
        RECT  6.375 0.275 8.000 0.365 ;
        RECT  6.370 1.435 8.000 1.525 ;
        RECT  7.100 0.780 7.250 0.890 ;
        RECT  7.000 0.505 7.100 1.315 ;
        RECT  6.565 0.505 7.000 0.615 ;
        RECT  6.735 1.205 7.000 1.315 ;
        RECT  6.765 0.750 6.875 1.095 ;
        RECT  6.585 1.005 6.765 1.095 ;
        RECT  6.495 1.005 6.585 1.320 ;
        RECT  6.475 0.505 6.565 0.890 ;
        RECT  5.985 1.230 6.495 1.320 ;
        RECT  6.390 0.780 6.475 0.890 ;
        RECT  6.275 0.275 6.375 0.645 ;
        RECT  6.200 1.410 6.370 1.525 ;
        RECT  6.185 0.970 6.280 1.140 ;
        RECT  5.780 1.435 6.200 1.525 ;
        RECT  6.095 0.275 6.185 1.140 ;
        RECT  5.935 0.275 6.095 0.365 ;
        RECT  5.985 0.475 6.005 0.645 ;
        RECT  5.895 0.475 5.985 1.320 ;
        RECT  5.765 0.255 5.935 0.365 ;
        RECT  5.715 0.455 5.805 1.155 ;
        RECT  5.690 1.265 5.780 1.525 ;
        RECT  5.200 0.275 5.765 0.365 ;
        RECT  5.655 0.455 5.715 0.645 ;
        RECT  5.380 1.045 5.715 1.155 ;
        RECT  4.650 1.265 5.690 1.355 ;
        RECT  5.560 0.735 5.625 0.905 ;
        RECT  5.470 0.475 5.560 0.905 ;
        RECT  5.145 0.475 5.470 0.565 ;
        RECT  5.280 0.735 5.380 1.155 ;
        RECT  5.030 0.255 5.200 0.365 ;
        RECT  5.055 0.475 5.145 1.175 ;
        RECT  4.915 0.475 5.055 0.575 ;
        RECT  4.865 1.065 5.055 1.175 ;
        RECT  4.815 0.275 5.030 0.365 ;
        RECT  4.775 0.765 4.930 0.875 ;
        RECT  4.725 0.275 4.815 0.675 ;
        RECT  4.685 0.765 4.775 1.175 ;
        RECT  4.595 0.585 4.725 0.675 ;
        RECT  4.470 1.085 4.685 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.485 0.585 4.595 0.925 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.350 0.585 4.485 0.675 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.290 0.280 4.350 0.995 ;
        RECT  4.255 0.280 4.290 1.165 ;
        RECT  4.220 0.280 4.255 0.470 ;
        RECT  4.180 0.905 4.255 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.685 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.215 0.275 3.440 0.415 ;
        RECT  3.330 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.330 1.345 ;
        RECT  3.220 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.220 0.610 ;
        RECT  2.610 1.045 3.220 1.135 ;
        RECT  1.700 0.275 3.215 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQNXD4

MACRO SEDFQXD0
    CLASS CORE ;
    FOREIGN SEDFQXD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.295 7.350 1.490 ;
        RECT  7.215 0.295 7.250 0.465 ;
        RECT  7.215 1.280 7.250 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0724 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 7.400 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.485 1.635 7.400 1.965 ;
        RECT  5.315 1.445 5.485 1.965 ;
        RECT  4.930 1.635 5.315 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.035 0.275 7.125 1.525 ;
        RECT  6.340 0.275 7.035 0.365 ;
        RECT  6.335 1.435 7.035 1.525 ;
        RECT  6.855 0.505 6.945 1.290 ;
        RECT  6.565 0.505 6.855 0.615 ;
        RECT  6.705 1.180 6.855 1.290 ;
        RECT  6.655 0.750 6.765 1.090 ;
        RECT  6.570 1.000 6.655 1.090 ;
        RECT  6.480 1.000 6.570 1.305 ;
        RECT  6.475 0.505 6.565 0.890 ;
        RECT  5.950 1.215 6.480 1.305 ;
        RECT  6.355 0.780 6.475 0.890 ;
        RECT  6.240 0.275 6.340 0.645 ;
        RECT  6.165 1.395 6.335 1.525 ;
        RECT  6.150 0.955 6.245 1.125 ;
        RECT  5.745 1.435 6.165 1.525 ;
        RECT  6.060 0.275 6.150 1.125 ;
        RECT  5.900 0.275 6.060 0.365 ;
        RECT  5.950 0.475 5.970 0.645 ;
        RECT  5.860 0.475 5.950 1.305 ;
        RECT  5.730 0.255 5.900 0.365 ;
        RECT  5.680 0.455 5.770 1.155 ;
        RECT  5.655 1.265 5.745 1.525 ;
        RECT  5.165 0.275 5.730 0.365 ;
        RECT  5.620 0.455 5.680 0.645 ;
        RECT  5.345 1.045 5.680 1.155 ;
        RECT  4.650 1.265 5.655 1.355 ;
        RECT  5.525 0.735 5.590 0.905 ;
        RECT  5.435 0.475 5.525 0.905 ;
        RECT  5.155 0.475 5.435 0.565 ;
        RECT  5.245 0.735 5.345 1.155 ;
        RECT  4.995 0.255 5.165 0.365 ;
        RECT  5.065 0.475 5.155 1.175 ;
        RECT  4.880 0.475 5.065 0.575 ;
        RECT  4.875 1.065 5.065 1.175 ;
        RECT  4.780 0.275 4.995 0.365 ;
        RECT  4.785 0.765 4.940 0.875 ;
        RECT  4.695 0.765 4.785 1.175 ;
        RECT  4.690 0.275 4.780 0.675 ;
        RECT  4.470 1.085 4.695 1.175 ;
        RECT  4.600 0.585 4.690 0.675 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.490 0.585 4.600 0.925 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.350 0.585 4.490 0.675 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.290 0.280 4.350 0.995 ;
        RECT  4.255 0.280 4.290 1.165 ;
        RECT  4.230 0.280 4.255 0.470 ;
        RECT  4.180 0.905 4.255 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.685 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.215 0.275 3.440 0.415 ;
        RECT  3.330 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.330 1.345 ;
        RECT  3.220 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.220 0.610 ;
        RECT  2.610 1.045 3.220 1.135 ;
        RECT  1.700 0.275 3.215 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.315 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.315 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQXD0

MACRO SEDFQXD1
    CLASS CORE ;
    FOREIGN SEDFQXD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 0.295 7.350 1.490 ;
        RECT  7.215 0.295 7.250 0.665 ;
        RECT  7.215 1.050 7.250 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 7.400 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.485 1.635 7.400 1.965 ;
        RECT  5.315 1.445 5.485 1.965 ;
        RECT  4.930 1.635 5.315 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.035 0.275 7.125 1.525 ;
        RECT  6.340 0.275 7.035 0.365 ;
        RECT  6.335 1.435 7.035 1.525 ;
        RECT  6.855 0.505 6.945 1.290 ;
        RECT  6.565 0.505 6.855 0.615 ;
        RECT  6.705 1.180 6.855 1.290 ;
        RECT  6.655 0.750 6.765 1.090 ;
        RECT  6.570 1.000 6.655 1.090 ;
        RECT  6.480 1.000 6.570 1.305 ;
        RECT  6.475 0.505 6.565 0.890 ;
        RECT  5.950 1.215 6.480 1.305 ;
        RECT  6.355 0.780 6.475 0.890 ;
        RECT  6.240 0.275 6.340 0.645 ;
        RECT  6.165 1.395 6.335 1.525 ;
        RECT  6.150 0.955 6.245 1.125 ;
        RECT  5.745 1.435 6.165 1.525 ;
        RECT  6.060 0.275 6.150 1.125 ;
        RECT  5.900 0.275 6.060 0.365 ;
        RECT  5.950 0.475 5.970 0.645 ;
        RECT  5.860 0.475 5.950 1.305 ;
        RECT  5.730 0.255 5.900 0.365 ;
        RECT  5.680 0.455 5.770 1.155 ;
        RECT  5.655 1.265 5.745 1.525 ;
        RECT  5.165 0.275 5.730 0.365 ;
        RECT  5.620 0.455 5.680 0.645 ;
        RECT  5.345 1.045 5.680 1.155 ;
        RECT  4.650 1.265 5.655 1.355 ;
        RECT  5.525 0.735 5.590 0.905 ;
        RECT  5.435 0.475 5.525 0.905 ;
        RECT  5.155 0.475 5.435 0.565 ;
        RECT  5.245 0.735 5.345 1.155 ;
        RECT  4.995 0.255 5.165 0.365 ;
        RECT  5.065 0.475 5.155 1.175 ;
        RECT  4.880 0.475 5.065 0.575 ;
        RECT  4.875 1.065 5.065 1.175 ;
        RECT  4.780 0.275 4.995 0.365 ;
        RECT  4.785 0.765 4.940 0.875 ;
        RECT  4.695 0.765 4.785 1.175 ;
        RECT  4.690 0.275 4.780 0.675 ;
        RECT  4.470 1.085 4.695 1.175 ;
        RECT  4.600 0.585 4.690 0.675 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.490 0.585 4.600 0.925 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.350 0.585 4.490 0.675 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.290 0.280 4.350 0.995 ;
        RECT  4.255 0.280 4.290 1.165 ;
        RECT  4.230 0.280 4.255 0.470 ;
        RECT  4.180 0.905 4.255 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.685 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.215 0.275 3.440 0.415 ;
        RECT  3.330 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.330 1.345 ;
        RECT  3.220 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.220 0.610 ;
        RECT  2.610 1.045 3.220 1.135 ;
        RECT  1.700 0.275 3.215 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQXD1

MACRO SEDFQXD2
    CLASS CORE ;
    FOREIGN SEDFQXD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.150 0.475 7.275 0.645 ;
        RECT  7.150 1.130 7.275 1.300 ;
        RECT  7.050 0.475 7.150 1.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 7.600 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.445 1.635 7.600 1.965 ;
        RECT  5.275 1.445 5.445 1.965 ;
        RECT  4.930 1.635 5.275 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.385 0.275 7.475 1.525 ;
        RECT  6.300 0.275 7.385 0.365 ;
        RECT  6.295 1.435 7.385 1.525 ;
        RECT  6.870 0.505 6.960 1.270 ;
        RECT  6.530 0.505 6.870 0.615 ;
        RECT  6.655 1.160 6.870 1.270 ;
        RECT  6.670 0.750 6.780 1.070 ;
        RECT  6.530 0.980 6.670 1.070 ;
        RECT  6.440 0.505 6.530 0.890 ;
        RECT  6.440 0.980 6.530 1.305 ;
        RECT  6.315 0.780 6.440 0.890 ;
        RECT  5.910 1.205 6.440 1.305 ;
        RECT  6.200 0.275 6.300 0.645 ;
        RECT  6.125 1.395 6.295 1.525 ;
        RECT  6.110 1.005 6.245 1.115 ;
        RECT  5.705 1.435 6.125 1.525 ;
        RECT  6.020 0.275 6.110 1.115 ;
        RECT  5.860 0.275 6.020 0.365 ;
        RECT  5.910 0.475 5.930 0.645 ;
        RECT  5.820 0.475 5.910 1.305 ;
        RECT  5.690 0.255 5.860 0.365 ;
        RECT  5.640 0.455 5.730 1.155 ;
        RECT  5.615 1.265 5.705 1.525 ;
        RECT  5.125 0.275 5.690 0.365 ;
        RECT  5.580 0.455 5.640 0.645 ;
        RECT  5.310 1.045 5.640 1.155 ;
        RECT  4.650 1.265 5.615 1.355 ;
        RECT  5.490 0.735 5.550 0.905 ;
        RECT  5.400 0.475 5.490 0.905 ;
        RECT  5.105 0.475 5.400 0.565 ;
        RECT  5.210 0.735 5.310 1.155 ;
        RECT  4.955 0.255 5.125 0.365 ;
        RECT  5.015 0.475 5.105 1.175 ;
        RECT  4.840 0.475 5.015 0.575 ;
        RECT  4.845 1.065 5.015 1.175 ;
        RECT  4.555 0.275 4.955 0.365 ;
        RECT  4.755 0.695 4.910 0.805 ;
        RECT  4.665 0.695 4.755 1.175 ;
        RECT  4.470 1.085 4.665 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.445 0.275 4.555 0.995 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  4.300 0.275 4.445 0.365 ;
        RECT  4.290 0.905 4.445 0.995 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.190 0.275 4.300 0.490 ;
        RECT  4.180 0.905 4.290 1.165 ;
        RECT  4.080 0.625 4.185 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.650 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.175 0.275 3.440 0.415 ;
        RECT  3.290 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.290 1.345 ;
        RECT  3.180 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.180 0.610 ;
        RECT  2.610 1.045 3.180 1.135 ;
        RECT  1.700 0.275 3.175 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQXD2

MACRO SEDFQXD4
    CLASS CORE ;
    FOREIGN SEDFQXD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.250 0.295 8.350 0.665 ;
        RECT  8.250 1.070 8.350 1.440 ;
        RECT  7.950 0.295 8.250 1.440 ;
        RECT  7.665 0.295 7.950 0.665 ;
        RECT  7.665 1.070 7.950 1.440 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0493 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 8.600 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.030 1.635 8.600 1.965 ;
        RECT  5.860 1.445 6.030 1.965 ;
        RECT  5.460 1.635 5.860 1.965 ;
        RECT  5.290 1.445 5.460 1.965 ;
        RECT  4.930 1.635 5.290 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.665 0.295 7.850 0.665 ;
        RECT  7.665 1.070 7.850 1.440 ;
        RECT  7.475 0.275 7.565 1.525 ;
        RECT  6.785 0.275 7.475 0.365 ;
        RECT  6.790 1.435 7.475 1.525 ;
        RECT  7.295 0.505 7.385 1.315 ;
        RECT  6.975 0.505 7.295 0.615 ;
        RECT  7.145 1.205 7.295 1.315 ;
        RECT  7.095 0.750 7.205 1.115 ;
        RECT  7.015 1.025 7.095 1.115 ;
        RECT  6.925 1.025 7.015 1.305 ;
        RECT  6.885 0.505 6.975 0.890 ;
        RECT  6.415 1.215 6.925 1.305 ;
        RECT  6.800 0.780 6.885 0.890 ;
        RECT  6.620 1.395 6.790 1.525 ;
        RECT  6.685 0.275 6.785 0.645 ;
        RECT  6.595 0.955 6.690 1.125 ;
        RECT  6.235 1.435 6.620 1.525 ;
        RECT  6.505 0.275 6.595 1.125 ;
        RECT  6.345 0.275 6.505 0.365 ;
        RECT  6.325 0.475 6.415 1.305 ;
        RECT  6.175 0.255 6.345 0.365 ;
        RECT  6.145 0.455 6.235 1.175 ;
        RECT  6.145 1.265 6.235 1.525 ;
        RECT  5.155 0.275 6.175 0.365 ;
        RECT  5.700 0.455 6.145 0.565 ;
        RECT  5.330 1.065 6.145 1.175 ;
        RECT  4.650 1.265 6.145 1.355 ;
        RECT  5.510 0.765 5.765 0.875 ;
        RECT  5.600 0.455 5.700 0.645 ;
        RECT  5.420 0.455 5.510 0.875 ;
        RECT  5.135 0.455 5.420 0.555 ;
        RECT  5.230 0.735 5.330 1.175 ;
        RECT  4.985 0.255 5.155 0.365 ;
        RECT  5.045 0.455 5.135 1.175 ;
        RECT  4.865 0.455 5.045 0.565 ;
        RECT  4.865 1.065 5.045 1.175 ;
        RECT  4.775 0.275 4.985 0.365 ;
        RECT  4.775 0.765 4.930 0.875 ;
        RECT  4.685 0.275 4.775 0.675 ;
        RECT  4.685 0.765 4.775 1.175 ;
        RECT  4.595 0.585 4.685 0.675 ;
        RECT  4.470 1.085 4.685 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.485 0.585 4.595 0.925 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.350 0.585 4.485 0.675 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.290 0.280 4.350 0.995 ;
        RECT  4.255 0.280 4.290 1.165 ;
        RECT  4.180 0.280 4.255 0.470 ;
        RECT  4.180 0.905 4.255 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.640 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.550 0.975 3.560 1.165 ;
        RECT  3.440 0.275 3.550 1.165 ;
        RECT  3.165 0.275 3.440 0.415 ;
        RECT  3.280 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.280 1.345 ;
        RECT  3.170 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.170 0.610 ;
        RECT  2.610 1.045 3.170 1.135 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  1.700 0.275 3.165 0.365 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFQXD4

MACRO SEDFXD0
    CLASS CORE ;
    FOREIGN SEDFXD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0610 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.550 1.030 6.640 1.140 ;
        RECT  6.550 0.565 6.620 0.675 ;
        RECT  6.450 0.565 6.550 1.140 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.495 7.750 1.290 ;
        RECT  7.625 0.495 7.650 0.665 ;
        RECT  7.625 1.060 7.650 1.290 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0724 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0220 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 7.800 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.510 1.635 7.800 1.965 ;
        RECT  7.340 1.505 7.510 1.965 ;
        RECT  5.500 1.635 7.340 1.965 ;
        RECT  5.330 1.445 5.500 1.965 ;
        RECT  4.930 1.635 5.330 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.445 0.305 7.535 1.410 ;
        RECT  7.055 0.305 7.445 0.415 ;
        RECT  7.205 1.320 7.445 1.410 ;
        RECT  7.265 0.565 7.355 1.185 ;
        RECT  6.970 0.565 7.265 0.675 ;
        RECT  7.005 1.075 7.265 1.185 ;
        RECT  7.095 1.320 7.205 1.525 ;
        RECT  7.065 0.770 7.175 0.965 ;
        RECT  6.825 0.875 7.065 0.965 ;
        RECT  6.735 0.305 7.055 0.400 ;
        RECT  6.915 1.075 7.005 1.525 ;
        RECT  5.760 1.435 6.915 1.525 ;
        RECT  6.735 0.875 6.825 1.325 ;
        RECT  6.545 0.305 6.735 0.425 ;
        RECT  5.965 1.235 6.735 1.325 ;
        RECT  6.165 1.055 6.280 1.145 ;
        RECT  6.075 0.275 6.165 1.145 ;
        RECT  5.915 0.275 6.075 0.365 ;
        RECT  5.965 0.475 5.985 0.645 ;
        RECT  5.875 0.475 5.965 1.325 ;
        RECT  5.745 0.255 5.915 0.365 ;
        RECT  5.695 0.455 5.785 1.155 ;
        RECT  5.670 1.265 5.760 1.525 ;
        RECT  5.180 0.275 5.745 0.365 ;
        RECT  5.635 0.455 5.695 0.645 ;
        RECT  5.360 1.045 5.695 1.155 ;
        RECT  4.650 1.265 5.670 1.355 ;
        RECT  5.540 0.735 5.605 0.905 ;
        RECT  5.450 0.475 5.540 0.905 ;
        RECT  5.155 0.475 5.450 0.565 ;
        RECT  5.260 0.735 5.360 1.155 ;
        RECT  5.010 0.255 5.180 0.365 ;
        RECT  5.065 0.475 5.155 1.175 ;
        RECT  4.895 0.475 5.065 0.575 ;
        RECT  4.875 1.065 5.065 1.175 ;
        RECT  4.795 0.275 5.010 0.365 ;
        RECT  4.785 0.765 4.940 0.875 ;
        RECT  4.705 0.275 4.795 0.630 ;
        RECT  4.695 0.765 4.785 1.175 ;
        RECT  4.600 0.540 4.705 0.630 ;
        RECT  4.470 1.085 4.695 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.490 0.540 4.600 0.925 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.350 0.540 4.490 0.630 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.290 0.280 4.350 0.995 ;
        RECT  4.255 0.280 4.290 1.165 ;
        RECT  4.240 0.280 4.255 0.470 ;
        RECT  4.180 0.905 4.255 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.695 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.225 0.275 3.440 0.415 ;
        RECT  3.340 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.340 1.345 ;
        RECT  3.230 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.230 0.610 ;
        RECT  2.610 1.045 3.230 1.135 ;
        RECT  1.700 0.275 3.225 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFXD0

MACRO SEDFXD1
    CLASS CORE ;
    FOREIGN SEDFXD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.505 7.550 1.170 ;
        RECT  7.285 0.505 7.450 0.615 ;
        RECT  7.425 1.070 7.450 1.170 ;
        RECT  7.315 1.070 7.425 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 0.295 7.950 1.490 ;
        RECT  7.825 0.295 7.850 0.665 ;
        RECT  7.815 1.070 7.850 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.590 -0.165 8.000 0.165 ;
        RECT  4.480 -0.165 4.590 0.490 ;
        RECT  1.310 -0.165 4.480 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.870 1.635 8.000 1.965 ;
        RECT  6.760 1.455 6.870 1.965 ;
        RECT  5.530 1.635 6.760 1.965 ;
        RECT  5.360 1.445 5.530 1.965 ;
        RECT  4.930 1.635 5.360 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.735 0.750 7.755 0.920 ;
        RECT  7.645 0.285 7.735 0.920 ;
        RECT  6.470 0.285 7.645 0.395 ;
        RECT  7.175 0.780 7.360 0.890 ;
        RECT  7.065 0.505 7.175 1.200 ;
        RECT  6.850 0.505 7.065 0.605 ;
        RECT  6.740 0.505 6.850 0.920 ;
        RECT  6.560 0.525 6.650 1.525 ;
        RECT  5.790 1.435 6.560 1.525 ;
        RECT  6.380 0.285 6.470 1.320 ;
        RECT  5.995 1.230 6.380 1.320 ;
        RECT  6.195 0.970 6.290 1.140 ;
        RECT  6.105 0.275 6.195 1.140 ;
        RECT  5.945 0.275 6.105 0.365 ;
        RECT  5.995 0.475 6.015 0.645 ;
        RECT  5.905 0.475 5.995 1.320 ;
        RECT  5.775 0.255 5.945 0.365 ;
        RECT  5.725 0.455 5.815 1.155 ;
        RECT  5.700 1.265 5.790 1.525 ;
        RECT  5.210 0.275 5.775 0.365 ;
        RECT  5.660 0.455 5.725 0.645 ;
        RECT  5.390 1.045 5.725 1.155 ;
        RECT  4.650 1.265 5.700 1.355 ;
        RECT  5.570 0.735 5.635 0.905 ;
        RECT  5.480 0.475 5.570 0.905 ;
        RECT  5.155 0.475 5.480 0.565 ;
        RECT  5.290 0.735 5.390 1.155 ;
        RECT  5.040 0.255 5.210 0.365 ;
        RECT  5.065 0.475 5.155 1.175 ;
        RECT  4.925 0.475 5.065 0.575 ;
        RECT  4.875 1.065 5.065 1.175 ;
        RECT  4.825 0.275 5.040 0.365 ;
        RECT  4.785 0.765 4.940 0.875 ;
        RECT  4.735 0.275 4.825 0.675 ;
        RECT  4.695 0.765 4.785 1.175 ;
        RECT  4.600 0.585 4.735 0.675 ;
        RECT  4.470 1.085 4.695 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.490 0.585 4.600 0.925 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.350 0.585 4.490 0.675 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.290 0.280 4.350 0.995 ;
        RECT  4.255 0.280 4.290 1.165 ;
        RECT  4.240 0.280 4.255 0.470 ;
        RECT  4.180 0.905 4.255 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.695 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.225 0.275 3.440 0.415 ;
        RECT  3.340 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.340 1.345 ;
        RECT  3.230 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.230 0.610 ;
        RECT  2.610 1.045 3.230 1.135 ;
        RECT  1.700 0.275 3.225 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFXD1

MACRO SEDFXD2
    CLASS CORE ;
    FOREIGN SEDFXD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.485 7.575 1.490 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 0.295 8.150 1.490 ;
        RECT  7.965 0.295 8.050 0.665 ;
        RECT  7.965 1.070 8.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 8.400 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.290 1.635 8.400 1.965 ;
        RECT  7.180 1.455 7.290 1.965 ;
        RECT  6.790 1.635 7.180 1.965 ;
        RECT  6.680 1.455 6.790 1.965 ;
        RECT  5.450 1.635 6.680 1.965 ;
        RECT  5.280 1.445 5.450 1.965 ;
        RECT  4.930 1.635 5.280 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.830 0.750 7.915 0.920 ;
        RECT  7.740 0.285 7.830 0.920 ;
        RECT  6.390 0.285 7.740 0.395 ;
        RECT  7.095 0.780 7.360 0.890 ;
        RECT  6.985 0.505 7.095 1.200 ;
        RECT  6.660 0.750 6.985 0.920 ;
        RECT  6.480 0.525 6.570 1.525 ;
        RECT  5.710 1.435 6.480 1.525 ;
        RECT  6.300 0.285 6.390 1.320 ;
        RECT  5.915 1.230 6.300 1.320 ;
        RECT  6.115 0.970 6.210 1.140 ;
        RECT  6.025 0.275 6.115 1.140 ;
        RECT  5.865 0.275 6.025 0.365 ;
        RECT  5.915 0.475 5.935 0.645 ;
        RECT  5.825 0.475 5.915 1.320 ;
        RECT  5.695 0.255 5.865 0.365 ;
        RECT  5.645 0.455 5.735 1.155 ;
        RECT  5.620 1.265 5.710 1.525 ;
        RECT  5.130 0.275 5.695 0.365 ;
        RECT  5.585 0.455 5.645 0.645 ;
        RECT  5.310 1.045 5.645 1.155 ;
        RECT  4.650 1.265 5.620 1.355 ;
        RECT  5.490 0.735 5.555 0.905 ;
        RECT  5.400 0.475 5.490 0.905 ;
        RECT  5.120 0.475 5.400 0.565 ;
        RECT  5.210 0.735 5.310 1.155 ;
        RECT  4.960 0.255 5.130 0.365 ;
        RECT  5.030 0.475 5.120 1.175 ;
        RECT  4.845 0.475 5.030 0.575 ;
        RECT  4.845 1.065 5.030 1.175 ;
        RECT  4.575 0.275 4.960 0.365 ;
        RECT  4.755 0.700 4.915 0.810 ;
        RECT  4.665 0.700 4.755 1.175 ;
        RECT  4.470 1.085 4.665 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.465 0.275 4.575 0.995 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  4.295 0.275 4.465 0.365 ;
        RECT  4.290 0.905 4.465 0.995 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.195 0.275 4.295 0.490 ;
        RECT  4.180 0.905 4.290 1.165 ;
        RECT  4.080 0.625 4.165 0.795 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.650 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.180 0.275 3.440 0.415 ;
        RECT  3.295 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.295 1.345 ;
        RECT  3.185 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.185 0.610 ;
        RECT  2.610 1.045 3.185 1.135 ;
        RECT  1.700 0.275 3.180 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFXD2

MACRO SEDFXD4
    CLASS CORE ;
    FOREIGN SEDFXD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0199 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.710 2.950 0.890 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.420 1.070 ;
        RECT  2.250 0.900 2.350 1.290 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.650 0.325 9.750 0.635 ;
        RECT  9.650 1.100 9.750 1.410 ;
        RECT  9.350 0.325 9.650 1.410 ;
        RECT  9.035 0.325 9.350 0.635 ;
        RECT  9.035 1.100 9.350 1.410 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.650 0.325 8.750 0.635 ;
        RECT  8.650 1.100 8.705 1.270 ;
        RECT  8.350 0.325 8.650 1.270 ;
        RECT  8.035 0.325 8.350 0.635 ;
        RECT  8.035 1.100 8.350 1.270 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0844 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.415 1.980 1.525 ;
        RECT  1.350 1.210 1.380 1.525 ;
        RECT  1.290 0.825 1.350 1.525 ;
        RECT  1.250 0.825 1.290 1.300 ;
        RECT  1.040 0.825 1.250 0.935 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.970 1.090 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0505 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.710 3.880 0.890 ;
        RECT  3.650 0.505 3.760 0.890 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.165 10.000 0.165 ;
        RECT  1.200 -0.165 1.310 0.440 ;
        RECT  0.000 -0.165 1.200 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.390 1.635 10.000 1.965 ;
        RECT  7.280 1.455 7.390 1.965 ;
        RECT  6.065 1.635 7.280 1.965 ;
        RECT  5.895 1.445 6.065 1.965 ;
        RECT  5.495 1.635 5.895 1.965 ;
        RECT  5.325 1.445 5.495 1.965 ;
        RECT  4.930 1.635 5.325 1.965 ;
        RECT  4.760 1.445 4.930 1.965 ;
        RECT  2.990 1.635 4.760 1.965 ;
        RECT  2.880 1.405 2.990 1.965 ;
        RECT  1.200 1.635 2.880 1.965 ;
        RECT  1.090 1.395 1.200 1.965 ;
        RECT  0.000 1.635 1.090 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.035 0.325 9.250 0.635 ;
        RECT  9.035 1.100 9.250 1.410 ;
        RECT  8.035 0.325 8.250 0.635 ;
        RECT  8.035 1.100 8.250 1.270 ;
        RECT  8.935 0.750 9.015 0.920 ;
        RECT  8.825 0.750 8.935 1.490 ;
        RECT  7.695 1.380 8.825 1.490 ;
        RECT  7.905 0.780 8.200 0.890 ;
        RECT  7.795 0.285 7.905 0.890 ;
        RECT  6.990 0.285 7.795 0.395 ;
        RECT  7.585 0.505 7.695 1.490 ;
        RECT  7.260 0.750 7.585 0.920 ;
        RECT  7.080 0.525 7.170 1.525 ;
        RECT  6.310 1.435 7.080 1.525 ;
        RECT  6.900 0.285 6.990 1.320 ;
        RECT  6.545 1.230 6.900 1.320 ;
        RECT  6.700 0.275 6.810 1.140 ;
        RECT  6.465 0.275 6.700 0.365 ;
        RECT  6.435 0.475 6.545 1.320 ;
        RECT  6.295 0.255 6.465 0.365 ;
        RECT  6.255 0.455 6.345 1.175 ;
        RECT  6.220 1.265 6.310 1.525 ;
        RECT  5.130 0.275 6.295 0.365 ;
        RECT  5.585 0.455 6.255 0.565 ;
        RECT  5.310 1.065 6.255 1.175 ;
        RECT  4.650 1.265 6.220 1.355 ;
        RECT  5.490 0.765 5.780 0.875 ;
        RECT  5.400 0.475 5.490 0.875 ;
        RECT  5.120 0.475 5.400 0.565 ;
        RECT  5.210 0.735 5.310 1.175 ;
        RECT  4.960 0.255 5.130 0.365 ;
        RECT  5.030 0.475 5.120 1.175 ;
        RECT  4.845 0.475 5.030 0.575 ;
        RECT  4.845 1.065 5.030 1.175 ;
        RECT  4.575 0.275 4.960 0.365 ;
        RECT  4.755 0.700 4.915 0.810 ;
        RECT  4.665 0.700 4.755 1.175 ;
        RECT  4.470 1.085 4.665 1.175 ;
        RECT  4.560 1.265 4.650 1.525 ;
        RECT  4.465 0.275 4.575 0.995 ;
        RECT  3.170 1.435 4.560 1.525 ;
        RECT  4.380 1.085 4.470 1.345 ;
        RECT  4.195 0.275 4.465 0.470 ;
        RECT  4.290 0.905 4.465 0.995 ;
        RECT  3.350 1.255 4.380 1.345 ;
        RECT  4.180 0.905 4.290 1.165 ;
        RECT  4.080 0.645 4.175 0.815 ;
        RECT  3.990 0.305 4.080 1.165 ;
        RECT  3.650 0.305 3.990 0.415 ;
        RECT  3.660 1.055 3.990 1.165 ;
        RECT  3.440 0.275 3.560 1.165 ;
        RECT  3.180 0.275 3.440 0.415 ;
        RECT  3.295 1.045 3.350 1.345 ;
        RECT  3.260 0.520 3.295 1.345 ;
        RECT  3.185 0.520 3.260 1.135 ;
        RECT  1.880 0.520 3.185 0.610 ;
        RECT  2.610 1.045 3.185 1.135 ;
        RECT  1.700 0.275 3.180 0.365 ;
        RECT  3.080 1.225 3.170 1.525 ;
        RECT  2.790 1.225 3.080 1.315 ;
        RECT  2.700 1.225 2.790 1.525 ;
        RECT  2.160 1.435 2.700 1.525 ;
        RECT  2.510 1.045 2.610 1.330 ;
        RECT  2.440 1.160 2.510 1.330 ;
        RECT  2.160 0.700 2.375 0.800 ;
        RECT  2.070 0.700 2.160 1.525 ;
        RECT  1.935 1.200 2.070 1.310 ;
        RECT  1.790 0.520 1.880 0.820 ;
        RECT  1.560 1.205 1.845 1.315 ;
        RECT  1.560 0.730 1.790 0.820 ;
        RECT  1.590 0.275 1.700 0.640 ;
        RECT  1.110 0.550 1.590 0.640 ;
        RECT  1.470 0.730 1.560 1.315 ;
        RECT  1.020 0.275 1.110 0.640 ;
        RECT  0.225 0.275 1.020 0.365 ;
        RECT  0.820 0.455 0.930 1.295 ;
        RECT  0.435 1.425 0.880 1.525 ;
        RECT  0.815 0.655 0.820 1.295 ;
        RECT  0.590 0.655 0.815 0.765 ;
        RECT  0.435 0.455 0.655 0.555 ;
        RECT  0.325 0.455 0.435 1.525 ;
        RECT  0.110 0.275 0.225 0.920 ;
    END
END SEDFXD4

MACRO TIEH
    CLASS CORE ;
    FOREIGN TIEH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.550 1.490 ;
        RECT  0.375 1.060 0.450 1.490 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 -0.165 0.600 0.165 ;
        RECT  0.115 -0.165 0.225 0.455 ;
        RECT  0.000 -0.165 0.115 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.635 0.600 1.965 ;
        RECT  0.115 1.050 0.225 1.965 ;
        RECT  0.000 1.635 0.115 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.375 0.275 0.485 0.665 ;
        RECT  0.310 0.565 0.375 0.665 ;
        RECT  0.200 0.565 0.310 0.940 ;
    END
END TIEH

MACRO TIEL
    CLASS CORE ;
    FOREIGN TIEL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.310 0.550 0.890 ;
        RECT  0.325 0.310 0.450 0.420 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 -0.165 0.600 0.165 ;
        RECT  0.115 -0.165 0.225 0.575 ;
        RECT  0.000 -0.165 0.115 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.635 0.600 1.965 ;
        RECT  0.115 1.280 0.225 1.965 ;
        RECT  0.000 1.635 0.115 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.375 1.070 0.485 1.480 ;
        RECT  0.310 1.070 0.375 1.170 ;
        RECT  0.200 0.730 0.310 1.170 ;
    END
END TIEL

MACRO XNR2D0
    CLASS CORE ;
    FOREIGN XNR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.510 1.950 1.330 ;
        RECT  1.755 0.510 1.850 0.620 ;
        RECT  1.755 1.220 1.850 1.330 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.555 0.910 ;
        RECT  1.375 0.740 1.450 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0565 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.640 -0.165 2.000 0.165 ;
        RECT  1.510 -0.165 1.640 0.420 ;
        RECT  0.375 -0.165 1.510 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.635 2.000 1.965 ;
        RECT  1.490 1.385 1.630 1.965 ;
        RECT  0.515 1.635 1.490 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.670 0.755 1.760 1.110 ;
        RECT  1.555 1.020 1.670 1.110 ;
        RECT  1.465 1.020 1.555 1.295 ;
        RECT  0.995 1.205 1.465 1.295 ;
        RECT  1.260 1.025 1.355 1.115 ;
        RECT  1.260 0.440 1.335 0.630 ;
        RECT  1.165 0.275 1.260 1.115 ;
        RECT  0.715 1.385 1.230 1.485 ;
        RECT  0.690 0.275 1.165 0.365 ;
        RECT  0.885 0.475 0.995 1.295 ;
        RECT  0.570 0.555 0.750 1.145 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.325 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.430 ;
        RECT  0.050 0.445 0.140 1.430 ;
    END
END XNR2D0

MACRO XNR2D1
    CLASS CORE ;
    FOREIGN XNR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.565 1.950 1.305 ;
        RECT  1.850 0.565 1.855 1.455 ;
        RECT  1.830 0.565 1.850 0.665 ;
        RECT  1.745 1.205 1.850 1.455 ;
        RECT  1.720 0.285 1.830 0.665 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.500 1.555 0.910 ;
        RECT  1.325 0.740 1.445 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0563 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.595 -0.165 2.000 0.165 ;
        RECT  1.400 -0.165 1.595 0.410 ;
        RECT  0.360 -0.165 1.400 0.165 ;
        RECT  0.360 0.510 0.475 0.620 ;
        RECT  0.270 -0.165 0.360 0.620 ;
        RECT  0.000 -0.165 0.270 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.635 2.000 1.965 ;
        RECT  1.430 1.415 1.600 1.965 ;
        RECT  0.475 1.635 1.430 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.655 0.775 1.755 1.110 ;
        RECT  1.615 1.020 1.655 1.110 ;
        RECT  1.525 1.020 1.615 1.305 ;
        RECT  0.975 1.205 1.525 1.305 ;
        RECT  1.220 1.015 1.330 1.115 ;
        RECT  1.220 0.315 1.290 0.425 ;
        RECT  1.120 0.315 1.220 1.115 ;
        RECT  0.750 1.415 1.165 1.525 ;
        RECT  0.470 0.315 1.120 0.415 ;
        RECT  0.865 0.505 0.975 1.305 ;
        RECT  0.670 0.530 0.770 1.125 ;
        RECT  0.660 1.215 0.750 1.525 ;
        RECT  0.575 0.530 0.670 0.640 ;
        RECT  0.570 1.015 0.670 1.125 ;
        RECT  0.185 1.215 0.660 1.305 ;
        RECT  0.140 1.215 0.185 1.450 ;
        RECT  0.140 0.445 0.180 0.615 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XNR2D1

MACRO XNR2D2
    CLASS CORE ;
    FOREIGN XNR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.565 1.950 1.305 ;
        RECT  1.850 0.565 1.855 1.455 ;
        RECT  1.830 0.565 1.850 0.665 ;
        RECT  1.745 1.205 1.850 1.455 ;
        RECT  1.720 0.285 1.830 0.665 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.500 1.555 0.910 ;
        RECT  1.325 0.740 1.445 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0563 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.090 -0.165 2.200 0.165 ;
        RECT  1.980 -0.165 2.090 0.475 ;
        RECT  1.570 -0.165 1.980 0.165 ;
        RECT  1.435 -0.165 1.570 0.410 ;
        RECT  0.360 -0.165 1.435 0.165 ;
        RECT  0.360 0.510 0.475 0.620 ;
        RECT  0.270 -0.165 0.360 0.620 ;
        RECT  0.000 -0.165 0.270 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.635 2.200 1.965 ;
        RECT  1.430 1.415 1.600 1.965 ;
        RECT  0.475 1.635 1.430 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.655 0.775 1.755 1.110 ;
        RECT  1.615 1.020 1.655 1.110 ;
        RECT  1.525 1.020 1.615 1.305 ;
        RECT  0.975 1.205 1.525 1.305 ;
        RECT  1.220 1.015 1.330 1.115 ;
        RECT  1.220 0.315 1.310 0.425 ;
        RECT  1.120 0.315 1.220 1.115 ;
        RECT  0.750 1.415 1.170 1.525 ;
        RECT  0.470 0.315 1.120 0.415 ;
        RECT  0.865 0.505 0.975 1.305 ;
        RECT  0.670 0.530 0.770 1.125 ;
        RECT  0.660 1.215 0.750 1.525 ;
        RECT  0.575 0.530 0.670 0.640 ;
        RECT  0.570 1.015 0.670 1.125 ;
        RECT  0.185 1.215 0.660 1.305 ;
        RECT  0.140 1.215 0.185 1.450 ;
        RECT  0.140 0.445 0.180 0.615 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XNR2D2

MACRO XNR2D4
    CLASS CORE ;
    FOREIGN XNR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.755 0.275 3.865 0.675 ;
        RECT  3.755 1.030 3.865 1.480 ;
        RECT  3.650 0.585 3.755 0.675 ;
        RECT  3.650 1.030 3.755 1.170 ;
        RECT  3.350 0.585 3.650 1.170 ;
        RECT  3.235 0.275 3.350 0.675 ;
        RECT  3.240 1.030 3.350 1.490 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1640 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.355 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1401 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.700 2.955 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.695 ;
        RECT  3.605 -0.165 4.015 0.165 ;
        RECT  3.495 -0.165 3.605 0.475 ;
        RECT  0.965 -0.165 3.495 0.165 ;
        RECT  0.855 -0.165 0.965 0.570 ;
        RECT  0.475 -0.165 0.855 0.165 ;
        RECT  0.305 -0.165 0.475 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.030 4.125 1.965 ;
        RECT  3.605 1.635 4.015 1.965 ;
        RECT  3.495 1.280 3.605 1.965 ;
        RECT  3.085 1.635 3.495 1.965 ;
        RECT  2.915 1.455 3.085 1.965 ;
        RECT  0.445 1.635 2.915 1.965 ;
        RECT  0.335 1.270 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.755 0.275 3.865 0.675 ;
        RECT  3.755 1.030 3.865 1.480 ;
        RECT  3.750 0.585 3.755 0.675 ;
        RECT  3.750 1.030 3.755 1.170 ;
        RECT  3.135 0.770 3.230 0.940 ;
        RECT  3.045 0.275 3.135 1.345 ;
        RECT  2.030 0.275 3.045 0.365 ;
        RECT  2.545 1.255 3.045 1.345 ;
        RECT  2.550 0.455 2.885 0.555 ;
        RECT  2.550 1.035 2.815 1.145 ;
        RECT  2.460 0.455 2.550 1.145 ;
        RECT  2.435 1.255 2.545 1.525 ;
        RECT  2.285 0.455 2.370 1.145 ;
        RECT  2.280 0.455 2.285 1.525 ;
        RECT  2.140 0.455 2.280 0.555 ;
        RECT  2.175 1.055 2.280 1.525 ;
        RECT  1.990 0.845 2.190 0.955 ;
        RECT  0.705 1.435 2.175 1.525 ;
        RECT  1.920 0.275 2.030 0.565 ;
        RECT  1.915 1.065 2.030 1.315 ;
        RECT  1.900 0.655 1.990 0.955 ;
        RECT  1.420 0.455 1.920 0.565 ;
        RECT  1.420 1.065 1.915 1.155 ;
        RECT  1.510 0.655 1.900 0.765 ;
        RECT  1.220 1.245 1.805 1.345 ;
        RECT  1.220 0.275 1.800 0.365 ;
        RECT  1.330 0.455 1.420 1.155 ;
        RECT  1.130 0.275 1.220 1.345 ;
        RECT  1.115 0.275 1.130 0.600 ;
        RECT  1.065 1.235 1.130 1.345 ;
        RECT  0.705 0.750 1.040 0.920 ;
        RECT  0.595 0.360 0.705 1.525 ;
        RECT  0.185 0.510 0.595 0.600 ;
        RECT  0.185 1.030 0.595 1.120 ;
        RECT  0.075 0.360 0.185 0.600 ;
        RECT  0.075 1.030 0.185 1.480 ;
    END
END XNR2D4

MACRO XNR3D0
    CLASS CORE ;
    FOREIGN XNR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.260 0.310 3.350 1.490 ;
        RECT  3.215 0.310 3.260 0.575 ;
        RECT  3.220 1.270 3.260 1.490 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.700 2.950 1.100 ;
        RECT  2.830 0.700 2.845 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0558 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.190 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0281 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.390 0.700 1.450 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.060 -0.165 3.400 0.165 ;
        RECT  2.950 -0.165 3.060 0.575 ;
        RECT  2.020 -0.165 2.950 0.165 ;
        RECT  1.925 -0.165 2.020 0.645 ;
        RECT  1.590 -0.165 1.925 0.165 ;
        RECT  1.460 -0.165 1.590 0.345 ;
        RECT  0.475 -0.165 1.460 0.165 ;
        RECT  0.305 -0.165 0.475 0.385 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 1.635 3.400 1.965 ;
        RECT  1.980 1.195 2.075 1.965 ;
        RECT  1.875 1.195 1.980 1.305 ;
        RECT  0.500 1.635 1.980 1.965 ;
        RECT  0.330 1.420 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 0.775 3.170 0.945 ;
        RECT  3.040 0.775 3.130 1.525 ;
        RECT  2.560 1.435 3.040 1.525 ;
        RECT  2.740 1.215 2.850 1.325 ;
        RECT  2.740 0.415 2.845 0.525 ;
        RECT  2.650 0.290 2.740 1.325 ;
        RECT  2.200 0.290 2.650 0.380 ;
        RECT  2.470 0.500 2.560 1.525 ;
        RECT  2.345 0.500 2.470 0.600 ;
        RECT  2.415 1.250 2.470 1.525 ;
        RECT  2.290 0.710 2.380 1.065 ;
        RECT  1.770 0.975 2.290 1.065 ;
        RECT  2.110 0.290 2.200 0.865 ;
        RECT  1.965 0.755 2.110 0.865 ;
        RECT  1.660 1.395 1.870 1.525 ;
        RECT  1.765 0.475 1.770 1.065 ;
        RECT  1.655 0.475 1.765 1.245 ;
        RECT  1.070 1.435 1.660 1.525 ;
        RECT  1.175 0.285 1.295 1.325 ;
        RECT  0.690 0.285 1.175 0.375 ;
        RECT  0.980 0.500 1.070 1.525 ;
        RECT  0.830 0.500 0.980 0.610 ;
        RECT  0.855 1.205 0.980 1.315 ;
        RECT  0.760 0.725 0.870 1.115 ;
        RECT  0.370 1.025 0.760 1.115 ;
        RECT  0.595 0.285 0.690 0.585 ;
        RECT  0.590 0.495 0.595 0.585 ;
        RECT  0.480 0.495 0.590 0.915 ;
        RECT  0.280 0.495 0.370 1.310 ;
        RECT  0.185 0.495 0.280 0.590 ;
        RECT  0.185 1.210 0.280 1.310 ;
        RECT  0.070 0.285 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.475 ;
    END
END XNR3D0

MACRO XNR3D1
    CLASS CORE ;
    FOREIGN XNR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.275 3.350 1.490 ;
        RECT  3.215 0.275 3.250 0.675 ;
        RECT  3.220 1.030 3.250 1.490 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.700 2.950 1.100 ;
        RECT  2.820 0.700 2.845 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0622 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.190 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.390 0.700 1.450 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.165 3.400 0.165 ;
        RECT  2.945 -0.165 3.070 0.575 ;
        RECT  2.010 -0.165 2.945 0.165 ;
        RECT  1.915 -0.165 2.010 0.645 ;
        RECT  1.550 -0.165 1.915 0.165 ;
        RECT  1.440 -0.165 1.550 0.345 ;
        RECT  0.475 -0.165 1.440 0.165 ;
        RECT  0.305 -0.165 0.475 0.385 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 1.635 3.400 1.965 ;
        RECT  1.980 1.195 2.075 1.965 ;
        RECT  1.875 1.195 1.980 1.305 ;
        RECT  0.500 1.635 1.980 1.965 ;
        RECT  0.330 1.420 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 0.750 3.160 0.920 ;
        RECT  3.040 0.750 3.130 1.515 ;
        RECT  2.550 1.425 3.040 1.515 ;
        RECT  2.730 1.215 2.850 1.325 ;
        RECT  2.730 0.415 2.835 0.525 ;
        RECT  2.640 0.290 2.730 1.325 ;
        RECT  2.190 0.290 2.640 0.380 ;
        RECT  2.460 0.490 2.550 1.515 ;
        RECT  2.335 0.490 2.460 0.600 ;
        RECT  2.415 1.250 2.460 1.515 ;
        RECT  2.280 0.710 2.370 1.065 ;
        RECT  1.765 0.975 2.280 1.065 ;
        RECT  2.100 0.290 2.190 0.865 ;
        RECT  1.965 0.755 2.100 0.865 ;
        RECT  1.660 1.395 1.870 1.525 ;
        RECT  1.760 0.975 1.765 1.245 ;
        RECT  1.655 0.475 1.760 1.245 ;
        RECT  1.070 1.435 1.660 1.525 ;
        RECT  1.165 0.285 1.275 1.325 ;
        RECT  0.690 0.285 1.165 0.375 ;
        RECT  0.980 0.500 1.070 1.525 ;
        RECT  0.800 0.500 0.980 0.610 ;
        RECT  0.855 1.230 0.980 1.340 ;
        RECT  0.760 0.725 0.870 1.125 ;
        RECT  0.370 1.035 0.760 1.125 ;
        RECT  0.595 0.285 0.690 0.585 ;
        RECT  0.590 0.495 0.595 0.585 ;
        RECT  0.480 0.495 0.590 0.915 ;
        RECT  0.280 0.495 0.370 1.310 ;
        RECT  0.185 0.495 0.280 0.590 ;
        RECT  0.185 1.220 0.280 1.310 ;
        RECT  0.070 0.285 0.185 0.590 ;
        RECT  0.075 1.220 0.185 1.475 ;
    END
END XNR3D1

MACRO XNR3D2
    CLASS CORE ;
    FOREIGN XNR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.365 4.350 1.140 ;
        RECT  3.905 0.365 4.250 0.475 ;
        RECT  4.065 1.040 4.250 1.140 ;
        RECT  3.955 1.040 4.065 1.470 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.795 3.750 1.300 ;
        RECT  3.555 0.795 3.650 0.965 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0545 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.480 1.555 0.890 ;
        RECT  1.330 0.760 1.445 0.890 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.080 -0.165 4.400 0.165 ;
        RECT  1.905 -0.165 2.080 0.600 ;
        RECT  1.570 -0.165 1.905 0.165 ;
        RECT  1.460 -0.165 1.570 0.335 ;
        RECT  0.365 -0.165 1.460 0.165 ;
        RECT  0.365 0.510 0.480 0.610 ;
        RECT  0.275 -0.165 0.365 0.610 ;
        RECT  0.000 -0.165 0.275 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 1.635 4.400 1.965 ;
        RECT  4.215 1.260 4.325 1.965 ;
        RECT  3.815 1.635 4.215 1.965 ;
        RECT  3.645 1.390 3.815 1.965 ;
        RECT  2.040 1.635 3.645 1.965 ;
        RECT  1.940 1.135 2.040 1.965 ;
        RECT  1.620 1.635 1.940 1.965 ;
        RECT  1.450 1.505 1.620 1.965 ;
        RECT  0.475 1.635 1.450 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.900 0.565 4.010 0.940 ;
        RECT  3.765 0.565 3.900 0.655 ;
        RECT  3.675 0.275 3.765 0.655 ;
        RECT  3.230 0.275 3.675 0.365 ;
        RECT  3.445 0.455 3.565 0.565 ;
        RECT  3.445 1.055 3.505 1.525 ;
        RECT  3.395 0.455 3.445 1.525 ;
        RECT  3.345 0.455 3.395 1.130 ;
        RECT  2.220 1.435 3.395 1.525 ;
        RECT  3.230 1.235 3.295 1.345 ;
        RECT  3.120 0.275 3.230 1.345 ;
        RECT  2.710 0.275 3.120 0.380 ;
        RECT  3.105 1.235 3.120 1.345 ;
        RECT  2.970 1.235 3.015 1.345 ;
        RECT  2.860 0.490 2.970 1.345 ;
        RECT  2.410 1.255 2.860 1.345 ;
        RECT  2.710 1.065 2.725 1.165 ;
        RECT  2.600 0.275 2.710 1.165 ;
        RECT  2.555 1.065 2.600 1.165 ;
        RECT  2.260 0.325 2.510 0.435 ;
        RECT  2.410 0.535 2.460 0.985 ;
        RECT  2.350 0.535 2.410 1.345 ;
        RECT  2.310 0.895 2.350 1.345 ;
        RECT  2.170 0.325 2.260 0.780 ;
        RECT  2.130 0.890 2.220 1.525 ;
        RECT  1.790 0.690 2.170 0.780 ;
        RECT  2.010 0.890 2.130 0.995 ;
        RECT  1.730 1.315 1.840 1.525 ;
        RECT  1.690 0.455 1.790 1.225 ;
        RECT  1.375 1.315 1.730 1.405 ;
        RECT  1.285 1.215 1.375 1.405 ;
        RECT  1.220 1.015 1.355 1.125 ;
        RECT  1.220 0.325 1.335 0.435 ;
        RECT  0.990 1.215 1.285 1.325 ;
        RECT  1.120 0.325 1.220 1.125 ;
        RECT  0.750 1.415 1.155 1.525 ;
        RECT  0.475 0.325 1.120 0.415 ;
        RECT  0.880 0.505 0.990 1.325 ;
        RECT  0.735 1.015 0.775 1.125 ;
        RECT  0.660 1.215 0.750 1.525 ;
        RECT  0.625 0.505 0.735 1.125 ;
        RECT  0.185 1.215 0.660 1.305 ;
        RECT  0.585 1.015 0.625 1.125 ;
        RECT  0.140 1.215 0.185 1.490 ;
        RECT  0.140 0.425 0.175 0.615 ;
        RECT  0.050 0.425 0.140 1.490 ;
    END
END XNR3D2

MACRO XNR3D4
    CLASS CORE ;
    FOREIGN XNR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.275 5.550 0.685 ;
        RECT  5.450 1.020 5.550 1.490 ;
        RECT  5.365 0.275 5.450 1.490 ;
        RECT  5.150 0.595 5.365 1.120 ;
        RECT  4.975 0.595 5.150 0.685 ;
        RECT  4.975 1.020 5.150 1.120 ;
        RECT  4.865 0.275 4.975 0.685 ;
        RECT  4.865 1.020 4.975 1.470 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.700 4.350 0.900 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0563 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.365 -0.165 5.800 0.165 ;
        RECT  0.365 0.510 0.480 0.610 ;
        RECT  0.275 -0.165 0.365 0.610 ;
        RECT  0.000 -0.165 0.275 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.635 5.800 1.965 ;
        RECT  2.990 1.415 3.160 1.965 ;
        RECT  0.475 1.635 2.990 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.975 0.595 5.050 0.685 ;
        RECT  4.975 1.020 5.050 1.120 ;
        RECT  4.865 0.275 4.975 0.685 ;
        RECT  4.865 1.020 4.975 1.470 ;
        RECT  4.725 0.780 5.000 0.890 ;
        RECT  4.635 0.310 4.725 1.410 ;
        RECT  3.720 0.310 4.635 0.400 ;
        RECT  3.715 1.320 4.635 1.410 ;
        RECT  3.905 0.500 4.525 0.610 ;
        RECT  3.905 1.085 4.525 1.195 ;
        RECT  3.815 0.500 3.905 1.195 ;
        RECT  2.890 0.815 3.815 0.905 ;
        RECT  3.630 0.310 3.720 0.455 ;
        RECT  3.615 0.995 3.715 1.410 ;
        RECT  3.425 0.615 3.655 0.725 ;
        RECT  3.115 0.345 3.630 0.455 ;
        RECT  3.125 0.995 3.615 1.085 ;
        RECT  3.425 1.175 3.525 1.525 ;
        RECT  3.255 0.545 3.425 0.725 ;
        RECT  3.230 1.175 3.425 1.285 ;
        RECT  2.780 0.635 3.255 0.725 ;
        RECT  3.035 0.995 3.125 1.315 ;
        RECT  3.025 0.345 3.115 0.545 ;
        RECT  2.390 1.225 3.035 1.315 ;
        RECT  2.545 0.455 3.025 0.545 ;
        RECT  2.685 1.025 2.895 1.135 ;
        RECT  2.285 0.275 2.870 0.365 ;
        RECT  2.690 0.635 2.780 0.830 ;
        RECT  1.850 1.435 2.720 1.525 ;
        RECT  2.390 0.720 2.690 0.830 ;
        RECT  2.300 1.025 2.685 1.115 ;
        RECT  2.435 0.455 2.545 0.630 ;
        RECT  2.285 1.025 2.300 1.315 ;
        RECT  2.190 0.275 2.285 1.315 ;
        RECT  2.175 0.275 2.190 1.125 ;
        RECT  1.220 1.015 1.850 1.125 ;
        RECT  1.760 1.215 1.850 1.525 ;
        RECT  1.220 0.325 1.835 0.435 ;
        RECT  0.985 1.215 1.760 1.325 ;
        RECT  1.120 0.325 1.220 1.125 ;
        RECT  0.750 1.415 1.150 1.525 ;
        RECT  0.475 0.325 1.120 0.415 ;
        RECT  0.875 0.505 0.985 1.325 ;
        RECT  0.735 1.015 0.775 1.125 ;
        RECT  0.660 1.215 0.750 1.525 ;
        RECT  0.625 0.505 0.735 1.125 ;
        RECT  0.185 1.215 0.660 1.305 ;
        RECT  0.570 1.015 0.625 1.125 ;
        RECT  0.140 1.215 0.185 1.490 ;
        RECT  0.140 0.425 0.175 0.615 ;
        RECT  0.050 0.425 0.140 1.490 ;
    END
END XNR3D4

MACRO XNR4D0
    CLASS CORE ;
    FOREIGN XNR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.510 3.350 1.115 ;
        RECT  3.085 0.510 3.250 0.620 ;
        RECT  3.085 1.015 3.250 1.115 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0278 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.700 3.580 0.920 ;
        RECT  3.445 0.700 3.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0559 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.700 4.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.645 -0.165 5.000 0.165 ;
        RECT  4.555 -0.165 4.645 0.590 ;
        RECT  2.070 -0.165 4.555 0.165 ;
        RECT  1.970 -0.165 2.070 0.670 ;
        RECT  1.560 -0.165 1.970 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.625 1.635 5.000 1.965 ;
        RECT  4.455 1.445 4.625 1.965 ;
        RECT  2.075 1.635 4.455 1.965 ;
        RECT  1.965 1.405 2.075 1.965 ;
        RECT  0.515 1.635 1.965 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.860 0.445 4.950 1.355 ;
        RECT  4.755 0.445 4.860 0.590 ;
        RECT  4.175 1.250 4.860 1.355 ;
        RECT  4.325 0.275 4.435 0.940 ;
        RECT  3.795 0.275 4.325 0.365 ;
        RECT  4.085 0.750 4.175 1.355 ;
        RECT  3.995 0.495 4.105 0.610 ;
        RECT  3.905 0.495 3.995 1.505 ;
        RECT  3.415 1.415 3.905 1.505 ;
        RECT  3.685 0.275 3.795 1.305 ;
        RECT  3.585 1.210 3.685 1.305 ;
        RECT  3.325 1.225 3.415 1.505 ;
        RECT  2.975 1.225 3.325 1.315 ;
        RECT  2.795 1.435 3.215 1.525 ;
        RECT  2.885 0.275 2.975 1.315 ;
        RECT  2.250 0.275 2.885 0.365 ;
        RECT  2.705 0.455 2.795 1.525 ;
        RECT  2.565 0.455 2.705 0.565 ;
        RECT  2.515 1.405 2.705 1.525 ;
        RECT  2.525 0.825 2.615 1.315 ;
        RECT  1.790 1.225 2.525 1.315 ;
        RECT  2.340 0.475 2.430 1.115 ;
        RECT  2.200 1.015 2.340 1.115 ;
        RECT  2.160 0.275 2.250 0.890 ;
        RECT  2.060 0.780 2.160 0.890 ;
        RECT  1.065 1.425 1.860 1.525 ;
        RECT  1.790 0.465 1.820 0.835 ;
        RECT  1.710 0.465 1.790 1.315 ;
        RECT  1.680 0.725 1.710 1.315 ;
        RECT  1.190 0.275 1.295 1.245 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.975 1.205 1.065 1.525 ;
        RECT  0.970 1.205 0.975 1.295 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.450 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XNR4D0

MACRO XNR4D1
    CLASS CORE ;
    FOREIGN XNR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.510 3.350 1.115 ;
        RECT  3.085 0.510 3.250 0.620 ;
        RECT  3.085 1.015 3.250 1.115 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.700 3.580 0.920 ;
        RECT  3.445 0.700 3.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0563 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.700 4.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.645 -0.165 5.000 0.165 ;
        RECT  4.555 -0.165 4.645 0.590 ;
        RECT  3.550 -0.165 4.555 0.165 ;
        RECT  3.380 -0.165 3.550 0.405 ;
        RECT  2.070 -0.165 3.380 0.165 ;
        RECT  1.970 -0.165 2.070 0.670 ;
        RECT  1.560 -0.165 1.970 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.625 1.635 5.000 1.965 ;
        RECT  4.455 1.445 4.625 1.965 ;
        RECT  2.075 1.635 4.455 1.965 ;
        RECT  1.965 1.405 2.075 1.965 ;
        RECT  0.515 1.635 1.965 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.860 0.445 4.950 1.355 ;
        RECT  4.755 0.445 4.860 0.590 ;
        RECT  4.175 1.250 4.860 1.355 ;
        RECT  4.325 0.275 4.435 0.940 ;
        RECT  3.795 0.275 4.325 0.365 ;
        RECT  4.085 0.750 4.175 1.355 ;
        RECT  3.995 0.470 4.105 0.585 ;
        RECT  3.905 0.470 3.995 1.505 ;
        RECT  3.415 1.415 3.905 1.505 ;
        RECT  3.685 0.275 3.795 1.305 ;
        RECT  3.585 1.210 3.685 1.305 ;
        RECT  3.325 1.225 3.415 1.505 ;
        RECT  2.995 1.225 3.325 1.315 ;
        RECT  2.795 1.435 3.130 1.525 ;
        RECT  2.885 0.275 2.995 1.315 ;
        RECT  2.250 0.275 2.885 0.365 ;
        RECT  2.705 0.455 2.795 1.525 ;
        RECT  2.565 0.455 2.705 0.565 ;
        RECT  2.515 1.405 2.705 1.525 ;
        RECT  2.525 0.825 2.615 1.315 ;
        RECT  1.790 1.225 2.525 1.315 ;
        RECT  2.340 0.475 2.430 1.115 ;
        RECT  2.200 1.015 2.340 1.115 ;
        RECT  2.160 0.275 2.250 0.890 ;
        RECT  2.060 0.780 2.160 0.890 ;
        RECT  1.075 1.425 1.860 1.525 ;
        RECT  1.790 0.470 1.820 0.835 ;
        RECT  1.710 0.470 1.790 1.315 ;
        RECT  1.680 0.725 1.710 1.315 ;
        RECT  1.190 0.275 1.295 1.295 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.985 1.205 1.075 1.525 ;
        RECT  0.970 1.205 0.985 1.295 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.450 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XNR4D1

MACRO XNR4D2
    CLASS CORE ;
    FOREIGN XNR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.495 0.475 3.550 1.140 ;
        RECT  3.450 0.475 3.495 1.480 ;
        RECT  3.335 0.475 3.450 0.585 ;
        RECT  3.385 1.030 3.450 1.480 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0550 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 0.710 3.840 0.920 ;
        RECT  3.650 0.710 3.750 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 0.700 5.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.035 -0.165 5.400 0.165 ;
        RECT  4.845 -0.165 5.035 0.355 ;
        RECT  2.070 -0.165 4.845 0.165 ;
        RECT  1.970 -0.165 2.070 0.670 ;
        RECT  1.560 -0.165 1.970 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.055 1.635 5.400 1.965 ;
        RECT  4.945 1.210 5.055 1.965 ;
        RECT  3.755 1.635 4.945 1.965 ;
        RECT  3.630 1.270 3.755 1.965 ;
        RECT  2.075 1.635 3.630 1.965 ;
        RECT  1.965 1.405 2.075 1.965 ;
        RECT  0.515 1.635 1.965 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.260 0.445 5.350 1.360 ;
        RECT  4.435 0.445 5.260 0.545 ;
        RECT  5.155 1.250 5.260 1.360 ;
        RECT  4.745 0.845 4.845 1.525 ;
        RECT  4.025 1.435 4.745 1.525 ;
        RECT  4.655 0.635 4.735 0.735 ;
        RECT  4.545 0.635 4.655 1.280 ;
        RECT  4.420 1.170 4.545 1.280 ;
        RECT  4.335 0.445 4.435 1.045 ;
        RECT  4.305 0.875 4.335 1.045 ;
        RECT  4.205 1.170 4.330 1.280 ;
        RECT  4.205 0.275 4.245 0.680 ;
        RECT  4.115 0.275 4.205 1.280 ;
        RECT  2.995 0.275 4.115 0.365 ;
        RECT  3.935 0.490 4.025 1.525 ;
        RECT  3.835 0.490 3.935 0.600 ;
        RECT  3.905 1.125 3.935 1.525 ;
        RECT  3.115 0.730 3.225 1.515 ;
        RECT  2.795 1.405 3.115 1.515 ;
        RECT  2.885 0.275 2.995 1.290 ;
        RECT  2.250 0.275 2.885 0.365 ;
        RECT  2.705 0.455 2.795 1.515 ;
        RECT  2.565 0.455 2.705 0.565 ;
        RECT  2.515 1.405 2.705 1.515 ;
        RECT  2.525 0.825 2.615 1.315 ;
        RECT  1.790 1.225 2.525 1.315 ;
        RECT  2.340 0.475 2.430 1.115 ;
        RECT  2.200 1.015 2.340 1.115 ;
        RECT  2.160 0.275 2.250 0.890 ;
        RECT  2.060 0.780 2.160 0.890 ;
        RECT  1.080 1.425 1.860 1.525 ;
        RECT  1.790 0.470 1.820 0.835 ;
        RECT  1.710 0.470 1.790 1.315 ;
        RECT  1.680 0.725 1.710 1.315 ;
        RECT  1.190 0.275 1.295 1.290 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.990 1.205 1.080 1.525 ;
        RECT  0.970 1.205 0.990 1.295 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.450 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XNR4D2

MACRO XNR4D4
    CLASS CORE ;
    FOREIGN XNR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.555 4.135 0.655 ;
        RECT  3.955 1.025 4.065 1.485 ;
        RECT  3.850 1.025 3.955 1.125 ;
        RECT  3.550 0.555 3.850 1.125 ;
        RECT  3.355 0.555 3.550 0.655 ;
        RECT  3.495 1.025 3.550 1.125 ;
        RECT  3.385 1.025 3.495 1.485 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.370 0.800 4.470 0.910 ;
        RECT  4.250 0.700 4.370 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.640 0.700 5.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.675 -0.165 6.000 0.165 ;
        RECT  5.485 -0.165 5.675 0.355 ;
        RECT  4.400 -0.165 5.485 0.165 ;
        RECT  4.230 -0.165 4.400 0.285 ;
        RECT  3.830 -0.165 4.230 0.165 ;
        RECT  3.660 -0.165 3.830 0.285 ;
        RECT  2.070 -0.165 3.660 0.165 ;
        RECT  1.970 -0.165 2.070 0.670 ;
        RECT  1.560 -0.165 1.970 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.655 1.635 6.000 1.965 ;
        RECT  5.555 1.210 5.655 1.965 ;
        RECT  4.350 1.635 5.555 1.965 ;
        RECT  4.240 1.210 4.350 1.965 ;
        RECT  3.780 1.635 4.240 1.965 ;
        RECT  3.670 1.275 3.780 1.965 ;
        RECT  2.075 1.635 3.670 1.965 ;
        RECT  1.965 1.405 2.075 1.965 ;
        RECT  0.515 1.635 1.965 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.950 0.555 4.135 0.655 ;
        RECT  3.955 1.025 4.065 1.485 ;
        RECT  3.950 1.025 3.955 1.125 ;
        RECT  3.355 0.555 3.450 0.655 ;
        RECT  3.385 1.025 3.450 1.485 ;
        RECT  5.860 0.445 5.950 1.360 ;
        RECT  5.085 0.445 5.860 0.545 ;
        RECT  5.755 1.250 5.860 1.360 ;
        RECT  5.365 0.845 5.465 1.500 ;
        RECT  5.275 0.635 5.375 0.735 ;
        RECT  4.685 1.390 5.365 1.500 ;
        RECT  5.185 0.635 5.275 1.280 ;
        RECT  5.055 1.170 5.185 1.280 ;
        RECT  4.995 0.445 5.085 1.045 ;
        RECT  4.955 0.875 4.995 1.045 ;
        RECT  4.865 1.170 4.965 1.280 ;
        RECT  4.865 0.375 4.905 0.675 ;
        RECT  4.775 0.375 4.865 1.280 ;
        RECT  2.995 0.375 4.775 0.465 ;
        RECT  4.595 0.555 4.685 1.500 ;
        RECT  4.515 0.555 4.595 0.660 ;
        RECT  4.535 1.125 4.595 1.500 ;
        RECT  3.245 0.780 3.325 0.890 ;
        RECT  3.135 0.780 3.245 1.515 ;
        RECT  2.795 1.405 3.135 1.515 ;
        RECT  2.885 0.275 2.995 1.290 ;
        RECT  2.250 0.275 2.885 0.365 ;
        RECT  2.705 0.455 2.795 1.515 ;
        RECT  2.565 0.455 2.705 0.565 ;
        RECT  2.515 1.405 2.705 1.515 ;
        RECT  2.525 0.825 2.615 1.315 ;
        RECT  1.790 1.225 2.525 1.315 ;
        RECT  2.340 0.475 2.430 1.115 ;
        RECT  2.200 1.015 2.340 1.115 ;
        RECT  2.160 0.275 2.250 0.890 ;
        RECT  2.060 0.780 2.160 0.890 ;
        RECT  1.065 1.425 1.860 1.525 ;
        RECT  1.790 0.470 1.820 0.835 ;
        RECT  1.710 0.470 1.790 1.315 ;
        RECT  1.680 0.725 1.710 1.315 ;
        RECT  1.190 0.275 1.295 1.305 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.975 1.205 1.065 1.525 ;
        RECT  0.970 1.205 0.975 1.295 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.450 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XNR4D4

MACRO XOR2D0
    CLASS CORE ;
    FOREIGN XOR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.510 1.950 1.330 ;
        RECT  1.755 0.510 1.850 0.620 ;
        RECT  1.755 1.220 1.850 1.330 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.555 0.910 ;
        RECT  1.375 0.740 1.450 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0563 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.165 2.000 0.165 ;
        RECT  1.520 -0.165 1.630 0.420 ;
        RECT  0.375 -0.165 1.520 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.635 2.000 1.965 ;
        RECT  1.520 1.385 1.630 1.965 ;
        RECT  0.515 1.635 1.520 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.670 0.775 1.760 1.110 ;
        RECT  1.555 1.020 1.670 1.110 ;
        RECT  1.465 1.020 1.555 1.295 ;
        RECT  0.960 1.205 1.465 1.295 ;
        RECT  1.260 1.025 1.355 1.115 ;
        RECT  1.260 0.275 1.335 0.630 ;
        RECT  1.245 0.275 1.260 1.115 ;
        RECT  0.690 0.275 1.245 0.365 ;
        RECT  1.165 0.540 1.245 1.115 ;
        RECT  0.960 0.455 1.075 0.635 ;
        RECT  0.870 0.455 0.960 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.570 0.555 0.750 1.145 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.325 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.430 ;
        RECT  0.050 0.445 0.140 1.430 ;
    END
END XOR2D0

MACRO XOR2D1
    CLASS CORE ;
    FOREIGN XOR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.275 1.950 1.490 ;
        RECT  1.765 0.275 1.850 0.665 ;
        RECT  1.765 1.220 1.850 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0546 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.480 1.555 0.910 ;
        RECT  1.375 0.740 1.450 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0679 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.635 -0.165 2.000 0.165 ;
        RECT  1.465 -0.165 1.635 0.385 ;
        RECT  0.375 -0.165 1.465 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.635 2.000 1.965 ;
        RECT  1.455 1.385 1.645 1.965 ;
        RECT  0.515 1.635 1.455 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.670 0.775 1.760 1.110 ;
        RECT  1.575 1.020 1.670 1.110 ;
        RECT  1.485 1.020 1.575 1.295 ;
        RECT  0.960 1.205 1.485 1.295 ;
        RECT  1.260 0.275 1.335 0.630 ;
        RECT  1.260 1.025 1.335 1.115 ;
        RECT  1.245 0.275 1.260 1.115 ;
        RECT  0.690 0.275 1.245 0.365 ;
        RECT  1.165 0.540 1.245 1.115 ;
        RECT  0.960 0.455 1.075 0.635 ;
        RECT  0.870 0.455 0.960 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.570 0.555 0.750 1.145 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.325 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.430 ;
        RECT  0.050 0.445 0.140 1.430 ;
    END
END XOR2D1

MACRO XOR2D2
    CLASS CORE ;
    FOREIGN XOR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.865 0.570 1.950 1.290 ;
        RECT  1.850 0.275 1.865 1.455 ;
        RECT  1.755 0.275 1.850 0.665 ;
        RECT  1.755 1.200 1.850 1.455 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0547 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.480 1.555 0.910 ;
        RECT  1.375 0.740 1.450 0.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0677 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 -0.165 2.200 0.165 ;
        RECT  2.015 -0.165 2.125 0.475 ;
        RECT  1.635 -0.165 2.015 0.165 ;
        RECT  1.465 -0.165 1.635 0.385 ;
        RECT  0.375 -0.165 1.465 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 1.635 2.200 1.965 ;
        RECT  2.025 1.345 2.125 1.965 ;
        RECT  1.630 1.635 2.025 1.965 ;
        RECT  1.440 1.385 1.630 1.965 ;
        RECT  0.475 1.635 1.440 1.965 ;
        RECT  0.305 1.395 0.475 1.965 ;
        RECT  0.000 1.635 0.305 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.670 0.775 1.760 1.090 ;
        RECT  1.575 1.000 1.670 1.090 ;
        RECT  1.485 1.000 1.575 1.295 ;
        RECT  0.980 1.205 1.485 1.295 ;
        RECT  1.260 1.025 1.370 1.115 ;
        RECT  1.260 0.275 1.340 0.630 ;
        RECT  1.235 0.275 1.260 1.115 ;
        RECT  0.690 0.275 1.235 0.365 ;
        RECT  1.165 0.540 1.235 1.115 ;
        RECT  0.980 0.455 1.075 0.635 ;
        RECT  0.890 0.455 0.980 1.295 ;
        RECT  0.735 1.385 0.885 1.485 ;
        RECT  0.680 0.545 0.780 1.115 ;
        RECT  0.645 1.205 0.735 1.485 ;
        RECT  0.600 0.275 0.690 0.420 ;
        RECT  0.570 0.545 0.680 0.655 ;
        RECT  0.590 1.015 0.680 1.115 ;
        RECT  0.175 1.205 0.645 1.295 ;
        RECT  0.475 0.315 0.600 0.420 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.205 0.175 1.430 ;
        RECT  0.050 0.445 0.140 1.430 ;
    END
END XOR2D2

MACRO XOR2D4
    CLASS CORE ;
    FOREIGN XOR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.275 3.870 0.675 ;
        RECT  3.760 1.030 3.870 1.480 ;
        RECT  3.650 0.585 3.760 0.675 ;
        RECT  3.650 1.030 3.760 1.170 ;
        RECT  3.355 0.585 3.650 1.170 ;
        RECT  3.350 0.275 3.355 1.170 ;
        RECT  3.240 0.275 3.350 0.675 ;
        RECT  3.245 1.030 3.350 1.490 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.1640 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.710 0.355 0.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1473 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.700 2.955 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.165 4.200 0.165 ;
        RECT  4.015 -0.165 4.125 0.695 ;
        RECT  3.605 -0.165 4.015 0.165 ;
        RECT  3.495 -0.165 3.605 0.475 ;
        RECT  0.965 -0.165 3.495 0.165 ;
        RECT  0.855 -0.165 0.965 0.570 ;
        RECT  0.475 -0.165 0.855 0.165 ;
        RECT  0.305 -0.165 0.475 0.405 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.635 4.200 1.965 ;
        RECT  4.015 1.030 4.125 1.965 ;
        RECT  3.605 1.635 4.015 1.965 ;
        RECT  3.495 1.280 3.605 1.965 ;
        RECT  3.085 1.635 3.495 1.965 ;
        RECT  2.915 1.455 3.085 1.965 ;
        RECT  0.445 1.635 2.915 1.965 ;
        RECT  0.335 1.270 0.445 1.965 ;
        RECT  0.000 1.635 0.335 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.760 0.275 3.870 0.675 ;
        RECT  3.760 1.030 3.870 1.480 ;
        RECT  3.750 0.585 3.760 0.675 ;
        RECT  3.750 1.030 3.760 1.170 ;
        RECT  3.135 0.770 3.230 0.940 ;
        RECT  3.045 0.275 3.135 1.345 ;
        RECT  2.030 0.275 3.045 0.365 ;
        RECT  2.545 1.255 3.045 1.345 ;
        RECT  2.550 0.455 2.885 0.565 ;
        RECT  2.550 1.035 2.815 1.145 ;
        RECT  2.460 0.455 2.550 1.145 ;
        RECT  2.435 1.255 2.545 1.525 ;
        RECT  2.285 0.455 2.370 1.145 ;
        RECT  2.280 0.455 2.285 1.525 ;
        RECT  2.140 0.455 2.280 0.555 ;
        RECT  2.175 1.055 2.280 1.525 ;
        RECT  1.990 0.845 2.190 0.955 ;
        RECT  0.705 1.435 2.175 1.525 ;
        RECT  1.920 0.275 2.030 0.565 ;
        RECT  1.915 1.065 2.030 1.315 ;
        RECT  1.900 0.655 1.990 0.955 ;
        RECT  1.420 0.455 1.920 0.565 ;
        RECT  1.420 1.065 1.915 1.155 ;
        RECT  1.510 0.655 1.900 0.765 ;
        RECT  1.220 1.245 1.805 1.345 ;
        RECT  1.220 0.275 1.800 0.365 ;
        RECT  1.330 0.455 1.420 1.155 ;
        RECT  1.130 0.275 1.220 1.345 ;
        RECT  1.115 0.275 1.130 0.600 ;
        RECT  1.065 1.235 1.130 1.345 ;
        RECT  0.705 0.750 1.040 0.920 ;
        RECT  0.595 0.360 0.705 1.525 ;
        RECT  0.185 0.510 0.595 0.600 ;
        RECT  0.185 1.030 0.595 1.120 ;
        RECT  0.075 0.360 0.185 0.600 ;
        RECT  0.075 1.030 0.185 1.480 ;
    END
END XOR2D4

MACRO XOR3D0
    CLASS CORE ;
    FOREIGN XOR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0760 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.260 0.310 3.350 1.490 ;
        RECT  3.215 0.310 3.260 0.575 ;
        RECT  3.220 1.270 3.260 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.700 2.950 1.100 ;
        RECT  2.830 0.700 2.845 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.190 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.390 0.700 1.450 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.060 -0.165 3.400 0.165 ;
        RECT  2.950 -0.165 3.060 0.575 ;
        RECT  2.020 -0.165 2.950 0.165 ;
        RECT  1.925 -0.165 2.020 0.645 ;
        RECT  1.580 -0.165 1.925 0.165 ;
        RECT  1.470 -0.165 1.580 0.345 ;
        RECT  0.475 -0.165 1.470 0.165 ;
        RECT  0.305 -0.165 0.475 0.385 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 1.635 3.400 1.965 ;
        RECT  1.980 1.195 2.075 1.965 ;
        RECT  1.875 1.195 1.980 1.305 ;
        RECT  0.500 1.635 1.980 1.965 ;
        RECT  0.330 1.420 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 0.775 3.170 0.945 ;
        RECT  3.040 0.775 3.130 1.525 ;
        RECT  2.560 1.435 3.040 1.525 ;
        RECT  2.740 1.215 2.850 1.325 ;
        RECT  2.740 0.415 2.845 0.525 ;
        RECT  2.650 0.290 2.740 1.325 ;
        RECT  2.200 0.290 2.650 0.380 ;
        RECT  2.470 0.500 2.560 1.525 ;
        RECT  2.345 0.500 2.470 0.600 ;
        RECT  2.415 1.250 2.470 1.525 ;
        RECT  2.290 0.710 2.380 1.065 ;
        RECT  1.770 0.975 2.290 1.065 ;
        RECT  2.110 0.290 2.200 0.865 ;
        RECT  1.965 0.755 2.110 0.865 ;
        RECT  1.660 1.395 1.870 1.525 ;
        RECT  1.765 0.475 1.770 1.065 ;
        RECT  1.655 0.475 1.765 1.245 ;
        RECT  1.070 1.435 1.660 1.525 ;
        RECT  1.175 0.285 1.295 1.325 ;
        RECT  0.690 0.285 1.175 0.375 ;
        RECT  0.980 0.500 1.070 1.525 ;
        RECT  0.875 0.500 0.980 0.610 ;
        RECT  0.855 1.205 0.980 1.315 ;
        RECT  0.760 0.795 0.870 1.115 ;
        RECT  0.370 1.025 0.760 1.115 ;
        RECT  0.595 0.285 0.690 0.585 ;
        RECT  0.590 0.495 0.595 0.585 ;
        RECT  0.480 0.495 0.590 0.915 ;
        RECT  0.280 0.495 0.370 1.310 ;
        RECT  0.185 0.495 0.280 0.590 ;
        RECT  0.185 1.210 0.280 1.310 ;
        RECT  0.070 0.285 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.475 ;
    END
END XOR3D0

MACRO XOR3D1
    CLASS CORE ;
    FOREIGN XOR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.260 0.275 3.350 1.490 ;
        RECT  3.215 0.275 3.260 0.690 ;
        RECT  3.220 1.030 3.260 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.700 2.950 1.100 ;
        RECT  2.830 0.700 2.845 0.920 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0564 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.700 0.190 0.920 ;
        RECT  0.050 0.700 0.150 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.390 0.700 1.450 0.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.060 -0.165 3.400 0.165 ;
        RECT  2.950 -0.165 3.060 0.575 ;
        RECT  2.020 -0.165 2.950 0.165 ;
        RECT  1.925 -0.165 2.020 0.645 ;
        RECT  1.580 -0.165 1.925 0.165 ;
        RECT  1.470 -0.165 1.580 0.345 ;
        RECT  0.475 -0.165 1.470 0.165 ;
        RECT  0.305 -0.165 0.475 0.385 ;
        RECT  0.000 -0.165 0.305 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 1.635 3.400 1.965 ;
        RECT  1.980 1.195 2.075 1.965 ;
        RECT  1.875 1.195 1.980 1.305 ;
        RECT  0.500 1.635 1.980 1.965 ;
        RECT  0.330 1.420 0.500 1.965 ;
        RECT  0.000 1.635 0.330 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 0.775 3.170 0.945 ;
        RECT  3.040 0.775 3.130 1.515 ;
        RECT  2.560 1.425 3.040 1.515 ;
        RECT  2.740 1.215 2.850 1.325 ;
        RECT  2.740 0.415 2.845 0.525 ;
        RECT  2.650 0.290 2.740 1.325 ;
        RECT  2.200 0.290 2.650 0.380 ;
        RECT  2.470 0.490 2.560 1.515 ;
        RECT  2.345 0.490 2.470 0.600 ;
        RECT  2.415 1.250 2.470 1.515 ;
        RECT  2.290 0.710 2.380 1.065 ;
        RECT  1.770 0.975 2.290 1.065 ;
        RECT  2.110 0.290 2.200 0.865 ;
        RECT  1.965 0.755 2.110 0.865 ;
        RECT  1.660 1.395 1.870 1.525 ;
        RECT  1.765 0.475 1.770 1.065 ;
        RECT  1.655 0.475 1.765 1.245 ;
        RECT  1.070 1.435 1.660 1.525 ;
        RECT  1.175 0.285 1.295 1.325 ;
        RECT  0.690 0.285 1.175 0.375 ;
        RECT  0.980 0.500 1.070 1.525 ;
        RECT  0.875 0.500 0.980 0.610 ;
        RECT  0.855 1.205 0.980 1.315 ;
        RECT  0.760 0.795 0.870 1.115 ;
        RECT  0.370 1.025 0.760 1.115 ;
        RECT  0.595 0.285 0.690 0.585 ;
        RECT  0.590 0.495 0.595 0.585 ;
        RECT  0.480 0.495 0.590 0.915 ;
        RECT  0.280 0.495 0.370 1.310 ;
        RECT  0.185 0.495 0.280 0.590 ;
        RECT  0.185 1.210 0.280 1.310 ;
        RECT  0.070 0.285 0.185 0.590 ;
        RECT  0.075 1.210 0.185 1.475 ;
    END
END XOR3D1

MACRO XOR3D2
    CLASS CORE ;
    FOREIGN XOR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.465 0.565 3.550 1.140 ;
        RECT  3.450 0.345 3.465 1.515 ;
        RECT  3.365 0.345 3.450 0.660 ;
        RECT  3.355 1.050 3.450 1.515 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 1.030 3.155 1.490 ;
        RECT  3.045 0.730 3.095 1.490 ;
        RECT  3.005 0.730 3.045 1.120 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.555 1.100 ;
        RECT  1.360 0.700 1.450 0.910 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.165 3.800 0.165 ;
        RECT  3.615 -0.165 3.725 0.465 ;
        RECT  2.105 -0.165 3.615 0.165 ;
        RECT  1.935 -0.165 2.105 0.355 ;
        RECT  1.620 -0.165 1.935 0.165 ;
        RECT  1.450 -0.165 1.620 0.345 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.525 0.500 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 1.635 3.800 1.965 ;
        RECT  3.615 1.255 3.725 1.965 ;
        RECT  2.040 1.635 3.615 1.965 ;
        RECT  1.940 1.130 2.040 1.965 ;
        RECT  1.620 1.635 1.940 1.965 ;
        RECT  1.450 1.515 1.620 1.965 ;
        RECT  0.515 1.635 1.450 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.275 0.770 3.345 0.940 ;
        RECT  3.185 0.275 3.275 0.940 ;
        RECT  2.665 0.275 3.185 0.365 ;
        RECT  2.915 0.465 3.000 0.575 ;
        RECT  2.915 1.230 2.955 1.525 ;
        RECT  2.825 0.465 2.915 1.525 ;
        RECT  2.795 0.465 2.825 0.575 ;
        RECT  2.220 1.435 2.825 1.525 ;
        RECT  2.665 1.155 2.690 1.345 ;
        RECT  2.555 0.275 2.665 1.345 ;
        RECT  2.325 0.275 2.435 0.535 ;
        RECT  2.320 0.625 2.430 1.345 ;
        RECT  1.790 0.445 2.325 0.535 ;
        RECT  2.170 0.625 2.320 0.725 ;
        RECT  2.130 0.850 2.220 1.525 ;
        RECT  2.030 0.850 2.130 0.960 ;
        RECT  1.730 1.315 1.840 1.525 ;
        RECT  1.680 0.445 1.790 1.225 ;
        RECT  1.285 1.315 1.730 1.405 ;
        RECT  1.255 1.015 1.340 1.115 ;
        RECT  1.255 0.275 1.300 0.595 ;
        RECT  1.195 1.205 1.285 1.405 ;
        RECT  1.160 0.275 1.255 1.115 ;
        RECT  0.970 1.205 1.195 1.295 ;
        RECT  0.690 0.275 1.160 0.365 ;
        RECT  0.970 0.455 1.070 0.565 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.860 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.185 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 1.260 0.185 1.470 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.050 0.445 0.140 1.470 ;
    END
END XOR3D2

MACRO XOR3D4
    CLASS CORE ;
    FOREIGN XOR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.275 5.550 0.685 ;
        RECT  5.450 1.020 5.550 1.490 ;
        RECT  5.365 0.275 5.450 1.490 ;
        RECT  5.150 0.595 5.365 1.120 ;
        RECT  4.975 0.595 5.150 0.685 ;
        RECT  4.975 1.020 5.150 1.120 ;
        RECT  4.865 0.275 4.975 0.685 ;
        RECT  4.850 1.020 4.975 1.490 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.700 4.350 0.900 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1658 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.750 0.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.375 -0.165 5.800 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.635 5.800 1.965 ;
        RECT  2.990 1.415 3.160 1.965 ;
        RECT  0.515 1.635 2.990 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.975 0.595 5.050 0.685 ;
        RECT  4.975 1.020 5.050 1.120 ;
        RECT  4.865 0.275 4.975 0.685 ;
        RECT  4.850 1.020 4.975 1.490 ;
        RECT  4.725 0.780 5.000 0.890 ;
        RECT  4.635 0.310 4.725 1.410 ;
        RECT  3.720 0.310 4.635 0.400 ;
        RECT  3.705 1.320 4.635 1.410 ;
        RECT  3.905 0.500 4.525 0.610 ;
        RECT  3.905 1.105 4.525 1.195 ;
        RECT  3.815 0.500 3.905 1.195 ;
        RECT  2.890 0.815 3.815 0.905 ;
        RECT  3.630 0.310 3.720 0.455 ;
        RECT  3.615 0.995 3.705 1.410 ;
        RECT  3.425 0.615 3.655 0.725 ;
        RECT  3.115 0.345 3.630 0.455 ;
        RECT  3.125 0.995 3.615 1.085 ;
        RECT  3.425 1.175 3.525 1.525 ;
        RECT  3.255 0.545 3.425 0.725 ;
        RECT  3.230 1.175 3.425 1.285 ;
        RECT  2.780 0.635 3.255 0.725 ;
        RECT  3.035 0.995 3.125 1.315 ;
        RECT  3.025 0.345 3.115 0.545 ;
        RECT  2.390 1.225 3.035 1.315 ;
        RECT  2.560 0.455 3.025 0.545 ;
        RECT  2.685 1.025 2.895 1.135 ;
        RECT  2.300 0.275 2.885 0.365 ;
        RECT  2.690 0.635 2.780 0.830 ;
        RECT  1.545 1.435 2.720 1.525 ;
        RECT  2.405 0.720 2.690 0.830 ;
        RECT  2.300 1.025 2.685 1.115 ;
        RECT  2.450 0.455 2.560 0.630 ;
        RECT  2.190 0.275 2.300 1.315 ;
        RECT  1.255 0.430 1.850 0.540 ;
        RECT  1.690 1.015 1.800 1.245 ;
        RECT  1.255 1.015 1.690 1.115 ;
        RECT  1.450 1.205 1.545 1.525 ;
        RECT  0.970 1.205 1.450 1.295 ;
        RECT  1.160 0.275 1.255 1.115 ;
        RECT  0.690 0.275 1.160 0.365 ;
        RECT  0.970 0.455 1.070 0.565 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.845 1.475 ;
        RECT  0.625 1.260 0.715 1.475 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.185 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 1.260 0.185 1.480 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.050 0.445 0.140 1.480 ;
    END
END XOR3D4

MACRO XOR4D0
    CLASS CORE ;
    FOREIGN XOR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.510 3.350 1.115 ;
        RECT  3.085 0.510 3.250 0.620 ;
        RECT  3.085 1.015 3.250 1.115 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0283 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.700 3.580 0.920 ;
        RECT  3.445 0.700 3.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0559 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.700 4.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.645 -0.165 5.000 0.165 ;
        RECT  4.555 -0.165 4.645 0.590 ;
        RECT  2.070 -0.165 4.555 0.165 ;
        RECT  1.970 -0.165 2.070 0.670 ;
        RECT  1.560 -0.165 1.970 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.625 1.635 5.000 1.965 ;
        RECT  4.455 1.445 4.625 1.965 ;
        RECT  2.075 1.635 4.455 1.965 ;
        RECT  1.965 1.405 2.075 1.965 ;
        RECT  0.515 1.635 1.965 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.860 0.445 4.950 1.355 ;
        RECT  4.755 0.445 4.860 0.590 ;
        RECT  4.175 1.250 4.860 1.355 ;
        RECT  4.325 0.275 4.435 0.940 ;
        RECT  3.795 0.275 4.325 0.365 ;
        RECT  4.085 0.750 4.175 1.355 ;
        RECT  3.995 0.495 4.105 0.610 ;
        RECT  3.905 0.495 3.995 1.525 ;
        RECT  3.415 1.435 3.905 1.525 ;
        RECT  3.685 0.275 3.795 1.305 ;
        RECT  3.585 1.210 3.685 1.305 ;
        RECT  3.325 1.225 3.415 1.525 ;
        RECT  2.985 1.225 3.325 1.315 ;
        RECT  2.795 1.435 3.215 1.525 ;
        RECT  2.885 0.275 2.985 1.315 ;
        RECT  2.250 0.275 2.885 0.365 ;
        RECT  2.705 0.500 2.795 1.525 ;
        RECT  2.540 0.500 2.705 0.610 ;
        RECT  2.515 1.405 2.705 1.525 ;
        RECT  2.525 0.825 2.615 1.315 ;
        RECT  1.790 1.225 2.525 1.315 ;
        RECT  2.340 0.475 2.430 1.115 ;
        RECT  2.200 1.015 2.340 1.115 ;
        RECT  2.160 0.275 2.250 0.890 ;
        RECT  2.060 0.780 2.160 0.890 ;
        RECT  1.065 1.425 1.860 1.525 ;
        RECT  1.790 0.465 1.820 0.835 ;
        RECT  1.710 0.465 1.790 1.315 ;
        RECT  1.680 0.725 1.710 1.315 ;
        RECT  1.190 0.275 1.295 1.220 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.975 1.205 1.065 1.525 ;
        RECT  0.970 1.205 0.975 1.295 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.450 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XOR4D0

MACRO XOR4D1
    CLASS CORE ;
    FOREIGN XOR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.510 3.350 1.115 ;
        RECT  3.085 0.510 3.250 0.620 ;
        RECT  3.085 1.015 3.250 1.115 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0655 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0548 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.700 3.580 0.920 ;
        RECT  3.445 0.700 3.550 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0653 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.640 0.700 4.750 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.645 -0.165 5.000 0.165 ;
        RECT  4.555 -0.165 4.645 0.590 ;
        RECT  3.550 -0.165 4.555 0.165 ;
        RECT  3.380 -0.165 3.550 0.405 ;
        RECT  2.070 -0.165 3.380 0.165 ;
        RECT  1.970 -0.165 2.070 0.670 ;
        RECT  1.560 -0.165 1.970 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.625 1.635 5.000 1.965 ;
        RECT  4.455 1.445 4.625 1.965 ;
        RECT  2.075 1.635 4.455 1.965 ;
        RECT  1.965 1.405 2.075 1.965 ;
        RECT  0.515 1.635 1.965 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.860 0.445 4.950 1.355 ;
        RECT  4.755 0.445 4.860 0.590 ;
        RECT  4.175 1.250 4.860 1.355 ;
        RECT  4.325 0.275 4.435 0.940 ;
        RECT  3.795 0.275 4.325 0.365 ;
        RECT  4.085 0.750 4.175 1.355 ;
        RECT  3.995 0.470 4.105 0.585 ;
        RECT  3.905 0.470 3.995 1.505 ;
        RECT  3.415 1.415 3.905 1.505 ;
        RECT  3.685 0.275 3.795 1.305 ;
        RECT  3.585 1.210 3.685 1.305 ;
        RECT  3.325 1.225 3.415 1.505 ;
        RECT  2.985 1.225 3.325 1.315 ;
        RECT  2.795 1.435 3.130 1.525 ;
        RECT  2.885 0.275 2.985 1.315 ;
        RECT  2.250 0.275 2.885 0.365 ;
        RECT  2.705 0.500 2.795 1.525 ;
        RECT  2.540 0.500 2.705 0.610 ;
        RECT  2.515 1.405 2.705 1.525 ;
        RECT  2.525 0.825 2.615 1.315 ;
        RECT  1.790 1.225 2.525 1.315 ;
        RECT  2.340 0.475 2.430 1.115 ;
        RECT  2.200 1.015 2.340 1.115 ;
        RECT  2.160 0.275 2.250 0.890 ;
        RECT  2.060 0.780 2.160 0.890 ;
        RECT  1.285 1.425 1.860 1.525 ;
        RECT  1.790 0.380 1.820 0.835 ;
        RECT  1.710 0.380 1.790 1.315 ;
        RECT  1.680 0.725 1.710 1.315 ;
        RECT  1.295 1.015 1.340 1.115 ;
        RECT  1.190 0.275 1.295 1.115 ;
        RECT  1.195 1.205 1.285 1.525 ;
        RECT  0.970 1.205 1.195 1.295 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  1.145 1.015 1.190 1.115 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.450 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XOR4D1

MACRO XOR4D2
    CLASS CORE ;
    FOREIGN XOR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.495 0.475 3.550 1.140 ;
        RECT  3.450 0.475 3.495 1.480 ;
        RECT  3.335 0.475 3.450 0.585 ;
        RECT  3.385 1.030 3.450 1.480 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0655 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.355 1.130 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 0.700 3.840 0.920 ;
        RECT  3.650 0.700 3.750 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0650 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 0.700 5.150 1.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.035 -0.165 5.400 0.165 ;
        RECT  4.845 -0.165 5.035 0.355 ;
        RECT  2.070 -0.165 4.845 0.165 ;
        RECT  1.970 -0.165 2.070 0.670 ;
        RECT  1.560 -0.165 1.970 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.055 1.635 5.400 1.965 ;
        RECT  4.945 1.210 5.055 1.965 ;
        RECT  3.755 1.635 4.945 1.965 ;
        RECT  3.630 1.270 3.755 1.965 ;
        RECT  2.075 1.635 3.630 1.965 ;
        RECT  1.965 1.405 2.075 1.965 ;
        RECT  0.515 1.635 1.965 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.260 0.445 5.350 1.360 ;
        RECT  4.435 0.445 5.260 0.545 ;
        RECT  5.155 1.250 5.260 1.360 ;
        RECT  4.745 0.845 4.845 1.525 ;
        RECT  4.025 1.435 4.745 1.525 ;
        RECT  4.655 0.635 4.735 0.735 ;
        RECT  4.545 0.635 4.655 1.280 ;
        RECT  4.420 1.170 4.545 1.280 ;
        RECT  4.335 0.445 4.435 1.045 ;
        RECT  4.305 0.875 4.335 1.045 ;
        RECT  4.205 1.170 4.330 1.280 ;
        RECT  4.205 0.275 4.245 0.635 ;
        RECT  4.115 0.275 4.205 1.280 ;
        RECT  2.985 0.275 4.115 0.365 ;
        RECT  3.935 0.475 4.025 1.525 ;
        RECT  3.835 0.475 3.935 0.585 ;
        RECT  3.905 1.125 3.935 1.525 ;
        RECT  3.115 0.730 3.225 1.515 ;
        RECT  2.795 1.405 3.115 1.515 ;
        RECT  2.885 0.275 2.985 1.290 ;
        RECT  2.250 0.275 2.885 0.365 ;
        RECT  2.705 0.500 2.795 1.515 ;
        RECT  2.540 0.500 2.705 0.610 ;
        RECT  2.515 1.405 2.705 1.515 ;
        RECT  2.525 0.825 2.615 1.315 ;
        RECT  1.790 1.225 2.525 1.315 ;
        RECT  2.340 0.475 2.430 1.115 ;
        RECT  2.200 1.015 2.340 1.115 ;
        RECT  2.160 0.275 2.250 0.890 ;
        RECT  2.060 0.780 2.160 0.890 ;
        RECT  1.285 1.425 1.860 1.525 ;
        RECT  1.790 0.380 1.820 0.835 ;
        RECT  1.710 0.380 1.790 1.315 ;
        RECT  1.680 0.725 1.710 1.315 ;
        RECT  1.295 1.015 1.340 1.115 ;
        RECT  1.190 0.275 1.295 1.115 ;
        RECT  1.195 1.205 1.285 1.525 ;
        RECT  0.970 1.205 1.195 1.295 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  1.145 1.015 1.190 1.115 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.175 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.140 1.260 0.175 1.450 ;
        RECT  0.050 0.445 0.140 1.450 ;
    END
END XOR4D2

MACRO XOR4D4
    CLASS CORE ;
    FOREIGN XOR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 1.800 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.515 4.260 0.625 ;
        RECT  4.100 1.040 4.210 1.470 ;
        RECT  4.050 1.040 4.100 1.135 ;
        RECT  3.750 0.515 4.050 1.135 ;
        RECT  3.530 0.515 3.750 0.625 ;
        RECT  3.690 1.040 3.750 1.135 ;
        RECT  3.580 1.040 3.690 1.470 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0655 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.710 0.365 1.100 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0553 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.700 1.550 1.100 ;
        RECT  1.385 0.700 1.450 0.910 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1105 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.845 0.700 4.955 1.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0651 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.450 0.700 6.550 1.100 ;
        RECT  6.390 0.700 6.450 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.285 -0.165 6.600 0.165 ;
        RECT  6.115 -0.165 6.285 0.385 ;
        RECT  1.560 -0.165 6.115 0.165 ;
        RECT  1.450 -0.165 1.560 0.590 ;
        RECT  0.375 -0.165 1.450 0.165 ;
        RECT  0.375 0.530 0.480 0.620 ;
        RECT  0.285 -0.165 0.375 0.620 ;
        RECT  0.000 -0.165 0.285 0.165 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.245 1.635 6.600 1.965 ;
        RECT  6.075 1.420 6.245 1.965 ;
        RECT  4.495 1.635 6.075 1.965 ;
        RECT  4.385 1.455 4.495 1.965 ;
        RECT  3.950 1.635 4.385 1.965 ;
        RECT  3.840 1.315 3.950 1.965 ;
        RECT  0.515 1.635 3.840 1.965 ;
        RECT  0.345 1.445 0.515 1.965 ;
        RECT  0.000 1.635 0.345 1.965 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.150 0.515 4.260 0.625 ;
        RECT  4.150 1.040 4.210 1.470 ;
        RECT  3.530 0.515 3.650 0.625 ;
        RECT  3.580 1.040 3.650 1.470 ;
        RECT  6.405 0.275 6.515 0.590 ;
        RECT  6.405 1.210 6.515 1.440 ;
        RECT  6.300 0.495 6.405 0.590 ;
        RECT  6.300 1.210 6.405 1.310 ;
        RECT  6.210 0.495 6.300 1.310 ;
        RECT  6.025 0.495 6.210 0.590 ;
        RECT  5.965 0.730 6.065 1.145 ;
        RECT  5.935 0.275 6.025 0.590 ;
        RECT  5.955 0.730 5.965 1.510 ;
        RECT  5.865 1.045 5.955 1.510 ;
        RECT  5.665 0.275 5.935 0.365 ;
        RECT  5.210 1.420 5.865 1.510 ;
        RECT  5.775 0.475 5.845 0.935 ;
        RECT  5.755 0.475 5.775 1.310 ;
        RECT  5.685 0.845 5.755 1.310 ;
        RECT  5.590 1.200 5.685 1.310 ;
        RECT  5.585 0.275 5.665 0.735 ;
        RECT  5.575 0.275 5.585 1.025 ;
        RECT  5.480 0.645 5.575 1.025 ;
        RECT  5.390 1.200 5.500 1.310 ;
        RECT  5.390 0.315 5.485 0.535 ;
        RECT  5.300 0.315 5.390 1.310 ;
        RECT  2.935 0.315 5.300 0.405 ;
        RECT  5.100 0.495 5.210 1.510 ;
        RECT  4.710 1.420 5.100 1.510 ;
        RECT  4.600 0.495 4.710 1.510 ;
        RECT  3.360 0.740 3.470 1.435 ;
        RECT  2.415 1.345 3.360 1.435 ;
        RECT  3.085 0.495 3.195 1.255 ;
        RECT  2.675 1.155 3.085 1.255 ;
        RECT  2.825 0.275 2.935 0.935 ;
        RECT  2.175 0.275 2.825 0.365 ;
        RECT  2.565 0.475 2.675 1.255 ;
        RECT  2.305 0.475 2.415 1.435 ;
        RECT  2.155 0.275 2.175 0.690 ;
        RECT  2.085 0.275 2.155 1.255 ;
        RECT  2.045 0.480 2.085 1.255 ;
        RECT  1.935 1.355 2.050 1.465 ;
        RECT  1.935 0.290 1.980 0.400 ;
        RECT  1.845 0.290 1.935 1.465 ;
        RECT  1.810 0.290 1.845 0.640 ;
        RECT  1.735 1.085 1.845 1.195 ;
        RECT  1.705 0.530 1.810 0.640 ;
        RECT  1.620 1.315 1.725 1.525 ;
        RECT  1.300 1.315 1.620 1.405 ;
        RECT  1.295 1.015 1.340 1.115 ;
        RECT  1.210 1.205 1.300 1.405 ;
        RECT  1.190 0.275 1.295 1.115 ;
        RECT  0.970 1.205 1.210 1.295 ;
        RECT  0.690 0.275 1.190 0.365 ;
        RECT  1.145 1.015 1.190 1.115 ;
        RECT  0.970 0.455 1.090 0.565 ;
        RECT  0.860 0.455 0.970 1.295 ;
        RECT  0.715 1.385 0.865 1.485 ;
        RECT  0.625 1.260 0.715 1.485 ;
        RECT  0.600 0.510 0.710 1.155 ;
        RECT  0.600 0.275 0.690 0.415 ;
        RECT  0.185 1.260 0.625 1.355 ;
        RECT  0.475 0.315 0.600 0.415 ;
        RECT  0.140 1.260 0.185 1.480 ;
        RECT  0.140 0.445 0.175 0.615 ;
        RECT  0.050 0.445 0.140 1.480 ;
    END
END XOR4D4

END LIBRARY
