module csa_tree_add1025_group_339_GENERIC_REAL(in_0, in_1, in_2, in_3,
     in_4, in_5, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( ( in_4 + in_5 )  + in_3 )  + in_2 )  + in_1 )  + in_0 )  ;"
  input [3:0] in_0, in_1, in_2, in_3, in_4, in_5;
  output [6:0] out_0;
  wire [3:0] in_0, in_1, in_2, in_3, in_4, in_5;
  wire [6:0] out_0;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_47, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_116, n_118, n_119, n_121, n_123, n_124, n_126;
  wire n_128, n_129, n_131, n_133, n_136, n_147, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_157, n_158;
  xor g1 (n_38, in_0[0], in_5[0]);
  and g15 (n_47, in_0[0], in_5[0]);
  xor g16 (n_62, in_4[0], in_1[0]);
  xor g2 (n_45, n_62, in_3[0]);
  nand g17 (n_63, in_4[0], in_1[0]);
  nand g18 (n_64, in_3[0], in_1[0]);
  nand g19 (n_65, in_4[0], in_3[0]);
  nand g20 (n_48, n_63, n_64, n_65);
  xor g21 (n_66, in_0[1], in_1[1]);
  xor g22 (n_49, n_66, in_3[1]);
  nand g3 (n_67, in_0[1], in_1[1]);
  nand g23 (n_68, in_3[1], in_1[1]);
  nand g24 (n_69, in_0[1], in_3[1]);
  nand g25 (n_52, n_67, n_68, n_69);
  xor g26 (n_70, in_5[1], in_4[1]);
  xor g27 (n_37, n_70, in_2[1]);
  nand g28 (n_71, in_5[1], in_4[1]);
  nand g4 (n_72, in_2[1], in_4[1]);
  nand g29 (n_73, in_5[1], in_2[1]);
  nand g30 (n_51, n_71, n_72, n_73);
  xor g31 (n_74, n_47, n_48);
  xor g32 (n_44, n_74, n_49);
  nand g33 (n_75, n_47, n_48);
  nand g34 (n_76, n_49, n_48);
  nand g5 (n_77, n_47, n_49);
  nand g35 (n_36, n_75, n_76, n_77);
  xor g36 (n_50, in_0[2], in_1[2]);
  and g37 (n_55, in_0[2], in_1[2]);
  xor g38 (n_78, in_3[2], in_4[2]);
  xor g39 (n_53, n_78, in_2[2]);
  nand g40 (n_79, in_3[2], in_4[2]);
  nand g41 (n_80, in_2[2], in_4[2]);
  nand g42 (n_81, in_3[2], in_2[2]);
  nand g6 (n_56, n_79, n_80, n_81);
  xor g43 (n_82, in_5[2], n_50);
  xor g44 (n_54, n_82, n_51);
  nand g45 (n_83, in_5[2], n_50);
  nand g46 (n_84, n_51, n_50);
  nand g47 (n_85, in_5[2], n_51);
  nand g48 (n_59, n_83, n_84, n_85);
  xor g49 (n_86, n_52, n_53);
  xor g50 (n_43, n_86, n_54);
  nand g51 (n_87, n_52, n_53);
  nand g52 (n_88, n_54, n_53);
  nand g53 (n_89, n_52, n_54);
  nand g54 (n_35, n_87, n_88, n_89);
  xor g55 (n_90, in_0[3], in_1[3]);
  xor g56 (n_57, n_90, in_3[3]);
  nand g57 (n_91, in_0[3], in_1[3]);
  nand g58 (n_92, in_3[3], in_1[3]);
  nand g59 (n_93, in_0[3], in_3[3]);
  nand g60 (n_61, n_91, n_92, n_93);
  xor g61 (n_94, in_4[3], in_2[3]);
  xor g62 (n_58, n_94, in_5[3]);
  nand g63 (n_95, in_4[3], in_2[3]);
  nand g64 (n_96, in_5[3], in_2[3]);
  nand g65 (n_97, in_4[3], in_5[3]);
  nand g66 (n_39, n_95, n_96, n_97);
  xor g67 (n_98, n_55, n_56);
  xor g68 (n_60, n_98, n_57);
  nand g69 (n_99, n_55, n_56);
  nand g70 (n_100, n_57, n_56);
  nand g71 (n_101, n_55, n_57);
  nand g72 (n_40, n_99, n_100, n_101);
  xor g73 (n_102, n_58, n_59);
  xor g74 (n_42, n_102, n_60);
  nand g75 (n_103, n_58, n_59);
  nand g76 (n_104, n_60, n_59);
  nand g77 (n_105, n_58, n_60);
  nand g78 (n_34, n_103, n_104, n_105);
  xor g79 (n_106, n_61, n_39);
  xor g80 (n_41, n_106, n_40);
  nand g81 (n_107, n_61, n_39);
  nand g82 (n_108, n_40, n_39);
  nand g83 (n_109, n_61, n_40);
  nand g84 (n_33, n_107, n_108, n_109);
  xor g85 (n_147, n_38, n_45);
  nand g86 (n_110, n_38, n_45);
  nand g87 (n_111, n_38, in_2[0]);
  nand g88 (n_112, n_45, in_2[0]);
  nand g89 (n_114, n_110, n_111, n_112);
  nor g90 (n_113, n_37, n_44);
  nand g7 (n_116, n_37, n_44);
  nor g8 (n_118, n_36, n_43);
  nand g9 (n_121, n_36, n_43);
  nor g10 (n_123, n_35, n_42);
  nand g11 (n_126, n_35, n_42);
  nor g12 (n_128, n_34, n_41);
  nand g13 (n_131, n_34, n_41);
  nand g96 (n_119, n_116, n_150);
  nand g99 (n_124, n_121, n_153);
  nand g102 (n_129, n_126, n_157);
  nand g105 (n_133, n_131, n_158);
  nand g107 (n_136, n_133, n_33);
  xnor g111 (out_0[1], n_114, n_151);
  xnor g113 (out_0[2], n_119, n_152);
  xnor g115 (out_0[3], n_124, n_154);
  xnor g117 (out_0[4], n_129, n_155);
  xor g122 (out_0[0], in_2[0], n_147);
  or g124 (n_150, n_113, wc);
  not gc (wc, n_114);
  or g125 (n_151, wc0, n_113);
  not gc0 (wc0, n_116);
  or g126 (n_152, wc1, n_118);
  not gc1 (wc1, n_121);
  or g127 (n_153, wc2, n_118);
  not gc2 (wc2, n_119);
  or g128 (n_154, wc3, n_123);
  not gc3 (wc3, n_126);
  or g129 (n_155, wc4, n_128);
  not gc4 (wc4, n_131);
  or g131 (n_157, wc5, n_123);
  not gc5 (wc5, n_124);
  or g132 (n_158, wc6, n_128);
  not gc6 (wc6, n_129);
  xor g133 (out_0[5], n_33, n_133);
  not g134 (out_0[6], n_136);
endmodule

module csa_tree_add1025_group_339_GENERIC(in_0, in_1, in_2, in_3, in_4,
     in_5, out_0);
  input [3:0] in_0, in_1, in_2, in_3, in_4, in_5;
  output [6:0] out_0;
  wire [3:0] in_0, in_1, in_2, in_3, in_4, in_5;
  wire [6:0] out_0;
  csa_tree_add1025_group_339_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .in_5 (in_5),
       .out_0 (out_0));
endmodule

module csa_tree_add_34_74_group_341_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( ( ( in_8 * in_9 )  + ( in_10 * in_11 )  )  + ( in_6 * in_7 )  )  + ( in_4 * in_5 )  )  + ( in_2 * in_3 )  )  + ( in_0 * in_1 )  )  ;"
  input [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  input [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  output [14:0] out_0;
  wire [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  wire [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  wire [14:0] out_0;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584;
  wire n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592;
  wire n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672;
  wire n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696;
  wire n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704;
  wire n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760;
  wire n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784;
  wire n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792;
  wire n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800;
  wire n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808;
  wire n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816;
  wire n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832;
  wire n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840;
  wire n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848;
  wire n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856;
  wire n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864;
  wire n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872;
  wire n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880;
  wire n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888;
  wire n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896;
  wire n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904;
  wire n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928;
  wire n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936;
  wire n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944;
  wire n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952;
  wire n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960;
  wire n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968;
  wire n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976;
  wire n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984;
  wire n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992;
  wire n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000;
  wire n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016;
  wire n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048;
  wire n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056;
  wire n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064;
  wire n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088;
  wire n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096;
  wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104;
  wire n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112;
  wire n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120;
  wire n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128;
  wire n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136;
  wire n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144;
  wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152;
  wire n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176;
  wire n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184;
  wire n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264;
  wire n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272;
  wire n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280;
  wire n_1281, n_1283, n_1285, n_1286, n_1288, n_1290, n_1291, n_1293;
  wire n_1295, n_1296, n_1298, n_1300, n_1301, n_1303, n_1305, n_1306;
  wire n_1308, n_1310, n_1311, n_1313, n_1315, n_1316, n_1318, n_1320;
  wire n_1321, n_1323, n_1325, n_1326, n_1328, n_1330, n_1331, n_1333;
  wire n_1335, n_1336, n_1338, n_1341, n_1344, n_1363, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1372, n_1373, n_1374, n_1375;
  wire n_1376, n_1377, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390;
  and g1 (n_119, in_0[0], in_1[0]);
  and g2 (n_124, in_0[1], in_1[0]);
  and g3 (n_142, in_0[2], in_1[0]);
  and g4 (n_173, in_0[3], in_1[0]);
  and g5 (n_223, in_0[4], in_1[0]);
  and g6 (n_282, in_0[5], in_1[0]);
  and g7 (n_345, in_0[6], in_1[0]);
  and g8 (n_410, in_0[7], in_1[0]);
  and g9 (n_125, in_0[0], in_1[1]);
  and g10 (n_143, in_0[1], in_1[1]);
  and g11 (n_174, in_0[2], in_1[1]);
  and g12 (n_224, in_0[3], in_1[1]);
  and g13 (n_283, in_0[4], in_1[1]);
  and g14 (n_346, in_0[5], in_1[1]);
  and g15 (n_411, in_0[6], in_1[1]);
  and g16 (n_476, in_0[7], in_1[1]);
  and g17 (n_151, in_0[0], in_1[2]);
  and g18 (n_189, in_0[1], in_1[2]);
  and g19 (n_239, in_0[2], in_1[2]);
  and g20 (n_298, in_0[3], in_1[2]);
  and g21 (n_361, in_0[4], in_1[2]);
  and g22 (n_426, in_0[5], in_1[2]);
  and g23 (n_477, in_0[6], in_1[2]);
  and g24 (n_533, in_0[7], in_1[2]);
  and g25 (n_175, in_0[0], in_1[3]);
  and g26 (n_225, in_0[1], in_1[3]);
  and g27 (n_284, in_0[2], in_1[3]);
  and g28 (n_347, in_0[3], in_1[3]);
  and g29 (n_412, in_0[4], in_1[3]);
  and g30 (n_487, in_0[5], in_1[3]);
  and g31 (n_534, in_0[6], in_1[3]);
  and g32 (n_577, in_0[7], in_1[3]);
  and g33 (n_122, in_2[0], in_3[0]);
  and g34 (n_133, in_2[1], in_3[0]);
  and g35 (n_144, in_2[2], in_3[0]);
  and g36 (n_182, in_2[3], in_3[0]);
  and g37 (n_232, in_2[4], in_3[0]);
  and g38 (n_291, in_2[5], in_3[0]);
  and g39 (n_354, in_2[6], in_3[0]);
  and g40 (n_419, in_2[7], in_3[0]);
  and g41 (n_126, in_2[0], in_3[1]);
  and g42 (n_104, in_2[1], in_3[1]);
  and g43 (n_190, in_2[2], in_3[1]);
  and g44 (n_240, in_2[3], in_3[1]);
  and g45 (n_299, in_2[4], in_3[1]);
  and g46 (n_362, in_2[5], in_3[1]);
  and g47 (n_427, in_2[6], in_3[1]);
  and g48 (n_478, in_2[7], in_3[1]);
  and g49 (n_152, in_2[0], in_3[2]);
  and g50 (n_194, in_2[1], in_3[2]);
  and g51 (n_244, in_2[2], in_3[2]);
  and g52 (n_303, in_2[3], in_3[2]);
  and g53 (n_366, in_2[4], in_3[2]);
  and g54 (n_431, in_2[5], in_3[2]);
  and g55 (n_484, in_2[6], in_3[2]);
  and g56 (n_541, in_2[7], in_3[2]);
  and g57 (n_176, in_2[0], in_3[3]);
  and g58 (n_226, in_2[1], in_3[3]);
  and g59 (n_285, in_2[2], in_3[3]);
  and g60 (n_348, in_2[3], in_3[3]);
  and g61 (n_413, in_2[4], in_3[3]);
  and g62 (n_488, in_2[5], in_3[3]);
  and g63 (n_535, in_2[6], in_3[3]);
  and g64 (n_578, in_2[7], in_3[3]);
  and g65 (n_118, in_4[0], in_5[0]);
  and g66 (n_132, in_4[1], in_5[0]);
  and g67 (n_157, in_4[2], in_5[0]);
  and g68 (n_179, in_4[3], in_5[0]);
  and g69 (n_229, in_4[4], in_5[0]);
  and g70 (n_288, in_4[5], in_5[0]);
  and g71 (n_351, in_4[6], in_5[0]);
  and g72 (n_416, in_4[7], in_5[0]);
  and g73 (n_134, in_4[0], in_5[1]);
  and g74 (n_145, in_4[1], in_5[1]);
  and g75 (n_183, in_4[2], in_5[1]);
  and g76 (n_233, in_4[3], in_5[1]);
  and g77 (n_292, in_4[4], in_5[1]);
  and g78 (n_355, in_4[5], in_5[1]);
  and g79 (n_420, in_4[6], in_5[1]);
  and g80 (n_491, in_4[7], in_5[1]);
  and g81 (n_148, in_4[0], in_5[2]);
  and g82 (n_186, in_4[1], in_5[2]);
  and g83 (n_236, in_4[2], in_5[2]);
  and g84 (n_295, in_4[3], in_5[2]);
  and g85 (n_358, in_4[4], in_5[2]);
  and g86 (n_423, in_4[5], in_5[2]);
  and g87 (n_479, in_4[6], in_5[2]);
  and g88 (n_538, in_4[7], in_5[2]);
  and g89 (n_191, in_4[0], in_5[3]);
  and g90 (n_241, in_4[1], in_5[3]);
  and g91 (n_300, in_4[2], in_5[3]);
  and g92 (n_363, in_4[3], in_5[3]);
  and g93 (n_428, in_4[4], in_5[3]);
  and g94 (n_482, in_4[5], in_5[3]);
  and g95 (n_542, in_4[6], in_5[3]);
  and g96 (n_581, in_4[7], in_5[3]);
  and g97 (n_123, in_6[0], in_7[0]);
  and g98 (n_135, in_6[1], in_7[0]);
  and g99 (n_149, in_6[2], in_7[0]);
  and g100 (n_193, in_6[3], in_7[0]);
  and g101 (n_243, in_6[4], in_7[0]);
  and g102 (n_302, in_6[5], in_7[0]);
  and g103 (n_365, in_6[6], in_7[0]);
  and g104 (n_430, in_6[7], in_7[0]);
  and g105 (n_128, in_6[0], in_7[1]);
  and g106 (n_150, in_6[1], in_7[1]);
  and g107 (n_195, in_6[2], in_7[1]);
  and g108 (n_245, in_6[3], in_7[1]);
  and g109 (n_304, in_6[4], in_7[1]);
  and g110 (n_367, in_6[5], in_7[1]);
  and g111 (n_432, in_6[6], in_7[1]);
  and g112 (n_485, in_6[7], in_7[1]);
  and g113 (n_153, in_6[0], in_7[2]);
  and g114 (n_196, in_6[1], in_7[2]);
  and g115 (n_246, in_6[2], in_7[2]);
  and g116 (n_305, in_6[3], in_7[2]);
  and g117 (n_368, in_6[4], in_7[2]);
  and g118 (n_433, in_6[5], in_7[2]);
  and g119 (n_486, in_6[6], in_7[2]);
  and g120 (n_544, in_6[7], in_7[2]);
  and g121 (n_177, in_6[0], in_7[3]);
  and g122 (n_227, in_6[1], in_7[3]);
  and g123 (n_286, in_6[2], in_7[3]);
  and g124 (n_349, in_6[3], in_7[3]);
  and g125 (n_414, in_6[4], in_7[3]);
  and g126 (n_489, in_6[5], in_7[3]);
  and g127 (n_536, in_6[6], in_7[3]);
  and g128 (n_579, in_6[7], in_7[3]);
  and g129 (n_121, in_8[0], in_9[0]);
  and g130 (n_131, in_8[1], in_9[0]);
  and g131 (n_156, in_8[2], in_9[0]);
  and g132 (n_178, in_8[3], in_9[0]);
  and g133 (n_228, in_8[4], in_9[0]);
  and g134 (n_287, in_8[5], in_9[0]);
  and g135 (n_350, in_8[6], in_9[0]);
  and g136 (n_415, in_8[7], in_9[0]);
  and g137 (n_130, in_8[0], in_9[1]);
  and g138 (n_155, in_8[1], in_9[1]);
  and g139 (n_180, in_8[2], in_9[1]);
  and g140 (n_230, in_8[3], in_9[1]);
  and g141 (n_289, in_8[4], in_9[1]);
  and g142 (n_352, in_8[5], in_9[1]);
  and g143 (n_417, in_8[6], in_9[1]);
  and g144 (n_490, in_8[7], in_9[1]);
  and g145 (n_154, in_8[0], in_9[2]);
  and g146 (n_181, in_8[1], in_9[2]);
  and g147 (n_231, in_8[2], in_9[2]);
  and g148 (n_290, in_8[3], in_9[2]);
  and g149 (n_353, in_8[4], in_9[2]);
  and g150 (n_418, in_8[5], in_9[2]);
  and g151 (n_492, in_8[6], in_9[2]);
  and g152 (n_537, in_8[7], in_9[2]);
  and g153 (n_184, in_8[0], in_9[3]);
  and g154 (n_234, in_8[1], in_9[3]);
  and g155 (n_293, in_8[2], in_9[3]);
  and g156 (n_356, in_8[3], in_9[3]);
  and g157 (n_421, in_8[4], in_9[3]);
  and g158 (n_493, in_8[5], in_9[3]);
  and g159 (n_539, in_8[6], in_9[3]);
  and g160 (n_580, in_8[7], in_9[3]);
  and g161 (n_120, in_10[0], in_11[0]);
  and g162 (n_129, in_10[1], in_11[0]);
  and g163 (n_146, in_10[2], in_11[0]);
  and g164 (n_185, in_10[3], in_11[0]);
  and g165 (n_235, in_10[4], in_11[0]);
  and g166 (n_294, in_10[5], in_11[0]);
  and g167 (n_357, in_10[6], in_11[0]);
  and g168 (n_422, in_10[7], in_11[0]);
  and g169 (n_127, in_10[0], in_11[1]);
  and g170 (n_147, in_10[1], in_11[1]);
  and g171 (n_187, in_10[2], in_11[1]);
  and g172 (n_237, in_10[3], in_11[1]);
  and g173 (n_296, in_10[4], in_11[1]);
  and g174 (n_359, in_10[5], in_11[1]);
  and g175 (n_424, in_10[6], in_11[1]);
  and g176 (n_480, in_10[7], in_11[1]);
  and g177 (n_103, in_10[0], in_11[2]);
  and g178 (n_188, in_10[1], in_11[2]);
  and g179 (n_238, in_10[2], in_11[2]);
  and g180 (n_297, in_10[3], in_11[2]);
  and g181 (n_360, in_10[4], in_11[2]);
  and g182 (n_425, in_10[5], in_11[2]);
  and g183 (n_481, in_10[6], in_11[2]);
  and g184 (n_540, in_10[7], in_11[2]);
  and g185 (n_192, in_10[0], in_11[3]);
  and g186 (n_242, in_10[1], in_11[3]);
  and g187 (n_301, in_10[2], in_11[3]);
  and g188 (n_364, in_10[3], in_11[3]);
  and g189 (n_429, in_10[4], in_11[3]);
  and g190 (n_483, in_10[5], in_11[3]);
  and g191 (n_543, in_10[6], in_11[3]);
  and g192 (n_582, in_10[7], in_11[3]);
  xor g363 (n_102, n_119, n_120);
  and g364 (n_136, n_119, n_120);
  xor g365 (n_621, n_121, n_122);
  xor g366 (n_117, n_621, n_123);
  nand g367 (n_622, n_121, n_122);
  nand g368 (n_623, n_123, n_122);
  nand g369 (n_624, n_121, n_123);
  nand g370 (n_137, n_622, n_623, n_624);
  xor g371 (n_625, n_124, n_125);
  xor g372 (n_139, n_625, n_126);
  nand g373 (n_626, n_124, n_125);
  nand g374 (n_627, n_126, n_125);
  nand g375 (n_628, n_124, n_126);
  nand g376 (n_161, n_626, n_627, n_628);
  xor g377 (n_629, n_127, n_128);
  xor g378 (n_138, n_629, n_129);
  nand g379 (n_630, n_127, n_128);
  nand g380 (n_631, n_129, n_128);
  nand g381 (n_632, n_127, n_129);
  nand g382 (n_158, n_630, n_631, n_632);
  xor g383 (n_633, n_130, n_131);
  xor g384 (n_141, n_633, n_132);
  nand g385 (n_634, n_130, n_131);
  nand g386 (n_635, n_132, n_131);
  nand g387 (n_636, n_130, n_132);
  nand g388 (n_160, n_634, n_635, n_636);
  xor g389 (n_637, n_133, n_134);
  xor g390 (n_140, n_637, n_135);
  nand g391 (n_638, n_133, n_134);
  nand g392 (n_639, n_135, n_134);
  nand g393 (n_640, n_133, n_135);
  nand g394 (n_159, n_638, n_639, n_640);
  xor g395 (n_641, n_136, n_137);
  xor g396 (n_101, n_641, n_138);
  nand g397 (n_642, n_136, n_137);
  nand g398 (n_643, n_138, n_137);
  nand g399 (n_644, n_136, n_138);
  nand g400 (n_169, n_642, n_643, n_644);
  xor g401 (n_645, n_139, n_140);
  xor g402 (n_116, n_645, n_141);
  nand g403 (n_646, n_139, n_140);
  nand g404 (n_647, n_141, n_140);
  nand g405 (n_648, n_139, n_141);
  nand g406 (n_168, n_646, n_647, n_648);
  xor g407 (n_649, n_142, n_143);
  xor g408 (n_164, n_649, n_144);
  nand g409 (n_650, n_142, n_143);
  nand g410 (n_651, n_144, n_143);
  nand g411 (n_652, n_142, n_144);
  nand g412 (n_202, n_650, n_651, n_652);
  xor g413 (n_653, n_145, n_146);
  xor g414 (n_162, n_653, n_147);
  nand g415 (n_654, n_145, n_146);
  nand g416 (n_655, n_147, n_146);
  nand g417 (n_656, n_145, n_147);
  nand g418 (n_198, n_654, n_655, n_656);
  xor g419 (n_657, n_148, n_103);
  xor g420 (n_163, n_657, n_104);
  nand g421 (n_658, n_148, n_103);
  nand g422 (n_659, n_104, n_103);
  nand g423 (n_660, n_148, n_104);
  nand g424 (n_200, n_658, n_659, n_660);
  xor g425 (n_661, n_149, n_150);
  xor g426 (n_165, n_661, n_151);
  nand g427 (n_662, n_149, n_150);
  nand g428 (n_663, n_151, n_150);
  nand g429 (n_664, n_149, n_151);
  nand g430 (n_203, n_662, n_663, n_664);
  xor g431 (n_665, n_152, n_153);
  xor g432 (n_166, n_665, n_154);
  nand g433 (n_666, n_152, n_153);
  nand g434 (n_667, n_154, n_153);
  nand g435 (n_668, n_152, n_154);
  nand g436 (n_199, n_666, n_667, n_668);
  xor g437 (n_669, n_155, n_156);
  xor g438 (n_167, n_669, n_157);
  nand g439 (n_670, n_155, n_156);
  nand g440 (n_671, n_157, n_156);
  nand g441 (n_672, n_155, n_157);
  nand g442 (n_201, n_670, n_671, n_672);
  xor g443 (n_673, n_158, n_159);
  xor g444 (n_170, n_673, n_160);
  nand g445 (n_674, n_158, n_159);
  nand g446 (n_675, n_160, n_159);
  nand g447 (n_676, n_158, n_160);
  nand g448 (n_211, n_674, n_675, n_676);
  xor g449 (n_677, n_161, n_162);
  xor g450 (n_172, n_677, n_163);
  nand g451 (n_678, n_161, n_162);
  nand g452 (n_679, n_163, n_162);
  nand g453 (n_680, n_161, n_163);
  nand g454 (n_215, n_678, n_679, n_680);
  xor g455 (n_681, n_164, n_165);
  xor g456 (n_171, n_681, n_166);
  nand g457 (n_682, n_164, n_165);
  nand g458 (n_683, n_166, n_165);
  nand g459 (n_684, n_164, n_166);
  nand g460 (n_214, n_682, n_683, n_684);
  xor g461 (n_685, n_167, n_168);
  xor g462 (n_100, n_685, n_169);
  nand g463 (n_686, n_167, n_168);
  nand g464 (n_687, n_169, n_168);
  nand g465 (n_688, n_167, n_169);
  nand g466 (n_220, n_686, n_687, n_688);
  xor g467 (n_689, n_170, n_171);
  xor g468 (n_115, n_689, n_172);
  nand g469 (n_690, n_170, n_171);
  nand g470 (n_691, n_172, n_171);
  nand g471 (n_692, n_170, n_172);
  nand g472 (n_221, n_690, n_691, n_692);
  xor g473 (n_197, n_173, n_174);
  and g474 (n_248, n_173, n_174);
  xor g475 (n_693, n_175, n_176);
  xor g476 (n_206, n_693, n_177);
  nand g477 (n_694, n_175, n_176);
  nand g478 (n_695, n_177, n_176);
  nand g479 (n_696, n_175, n_177);
  nand g480 (n_253, n_694, n_695, n_696);
  xor g481 (n_697, n_178, n_179);
  xor g482 (n_210, n_697, n_180);
  nand g483 (n_698, n_178, n_179);
  nand g484 (n_699, n_180, n_179);
  nand g485 (n_700, n_178, n_180);
  nand g486 (n_254, n_698, n_699, n_700);
  xor g487 (n_701, n_181, n_182);
  xor g488 (n_208, n_701, n_183);
  nand g489 (n_702, n_181, n_182);
  nand g490 (n_703, n_183, n_182);
  nand g491 (n_704, n_181, n_183);
  nand g492 (n_255, n_702, n_703, n_704);
  xor g493 (n_705, n_184, n_185);
  xor g494 (n_205, n_705, n_186);
  nand g495 (n_706, n_184, n_185);
  nand g496 (n_707, n_186, n_185);
  nand g497 (n_708, n_184, n_186);
  nand g498 (n_251, n_706, n_707, n_708);
  xor g499 (n_709, n_187, n_188);
  xor g500 (n_209, n_709, n_189);
  nand g501 (n_710, n_187, n_188);
  nand g502 (n_711, n_189, n_188);
  nand g503 (n_712, n_187, n_189);
  nand g504 (n_250, n_710, n_711, n_712);
  xor g505 (n_713, n_190, n_191);
  xor g506 (n_204, n_713, n_192);
  nand g507 (n_714, n_190, n_191);
  nand g508 (n_715, n_192, n_191);
  nand g509 (n_716, n_190, n_192);
  nand g510 (n_252, n_714, n_715, n_716);
  xor g511 (n_717, n_193, n_194);
  xor g512 (n_207, n_717, n_195);
  nand g513 (n_718, n_193, n_194);
  nand g514 (n_719, n_195, n_194);
  nand g515 (n_720, n_193, n_195);
  nand g516 (n_249, n_718, n_719, n_720);
  xor g517 (n_721, n_196, n_197);
  xor g518 (n_212, n_721, n_198);
  nand g519 (n_722, n_196, n_197);
  nand g520 (n_723, n_198, n_197);
  nand g521 (n_724, n_196, n_198);
  nand g522 (n_263, n_722, n_723, n_724);
  xor g523 (n_725, n_199, n_200);
  xor g524 (n_213, n_725, n_201);
  nand g525 (n_726, n_199, n_200);
  nand g526 (n_727, n_201, n_200);
  nand g527 (n_728, n_199, n_201);
  nand g528 (n_264, n_726, n_727, n_728);
  xor g529 (n_729, n_202, n_203);
  xor g530 (n_216, n_729, n_204);
  nand g531 (n_730, n_202, n_203);
  nand g532 (n_731, n_204, n_203);
  nand g533 (n_732, n_202, n_204);
  nand g534 (n_268, n_730, n_731, n_732);
  xor g535 (n_733, n_205, n_206);
  xor g536 (n_218, n_733, n_207);
  nand g537 (n_734, n_205, n_206);
  nand g538 (n_735, n_207, n_206);
  nand g539 (n_736, n_205, n_207);
  nand g540 (n_267, n_734, n_735, n_736);
  xor g541 (n_737, n_208, n_209);
  xor g542 (n_217, n_737, n_210);
  nand g543 (n_738, n_208, n_209);
  nand g544 (n_739, n_210, n_209);
  nand g545 (n_740, n_208, n_210);
  nand g546 (n_269, n_738, n_739, n_740);
  xor g547 (n_741, n_211, n_212);
  xor g548 (n_219, n_741, n_213);
  nand g549 (n_742, n_211, n_212);
  nand g550 (n_743, n_213, n_212);
  nand g551 (n_744, n_211, n_213);
  nand g552 (n_276, n_742, n_743, n_744);
  xor g553 (n_745, n_214, n_215);
  xor g554 (n_222, n_745, n_216);
  nand g555 (n_746, n_214, n_215);
  nand g556 (n_747, n_216, n_215);
  nand g557 (n_748, n_214, n_216);
  nand g558 (n_274, n_746, n_747, n_748);
  xor g559 (n_749, n_217, n_218);
  xor g560 (n_99, n_749, n_219);
  nand g561 (n_750, n_217, n_218);
  nand g562 (n_751, n_219, n_218);
  nand g563 (n_752, n_217, n_219);
  nand g564 (n_279, n_750, n_751, n_752);
  xor g565 (n_753, n_220, n_221);
  xor g566 (n_114, n_753, n_222);
  nand g567 (n_754, n_220, n_221);
  nand g568 (n_755, n_222, n_221);
  nand g569 (n_756, n_220, n_222);
  nand g570 (n_281, n_754, n_755, n_756);
  xor g571 (n_247, n_223, n_224);
  and g572 (n_306, n_223, n_224);
  xor g573 (n_757, n_225, n_226);
  xor g574 (n_261, n_757, n_227);
  nand g575 (n_758, n_225, n_226);
  nand g576 (n_759, n_227, n_226);
  nand g577 (n_760, n_225, n_227);
  nand g578 (n_309, n_758, n_759, n_760);
  xor g579 (n_761, n_228, n_229);
  xor g580 (n_258, n_761, n_230);
  nand g581 (n_762, n_228, n_229);
  nand g582 (n_763, n_230, n_229);
  nand g583 (n_764, n_228, n_230);
  nand g584 (n_310, n_762, n_763, n_764);
  xor g585 (n_765, n_231, n_232);
  xor g586 (n_260, n_765, n_233);
  nand g587 (n_766, n_231, n_232);
  nand g588 (n_767, n_233, n_232);
  nand g589 (n_768, n_231, n_233);
  nand g590 (n_312, n_766, n_767, n_768);
  xor g591 (n_769, n_234, n_235);
  xor g592 (n_259, n_769, n_236);
  nand g593 (n_770, n_234, n_235);
  nand g594 (n_771, n_236, n_235);
  nand g595 (n_772, n_234, n_236);
  nand g596 (n_308, n_770, n_771, n_772);
  xor g597 (n_773, n_237, n_238);
  xor g598 (n_256, n_773, n_239);
  nand g599 (n_774, n_237, n_238);
  nand g600 (n_775, n_239, n_238);
  nand g601 (n_776, n_237, n_239);
  nand g602 (n_313, n_774, n_775, n_776);
  xor g603 (n_777, n_240, n_241);
  xor g604 (n_262, n_777, n_242);
  nand g605 (n_778, n_240, n_241);
  nand g606 (n_779, n_242, n_241);
  nand g607 (n_780, n_240, n_242);
  nand g608 (n_311, n_778, n_779, n_780);
  xor g609 (n_781, n_243, n_244);
  xor g610 (n_257, n_781, n_245);
  nand g611 (n_782, n_243, n_244);
  nand g612 (n_783, n_245, n_244);
  nand g613 (n_784, n_243, n_245);
  nand g614 (n_307, n_782, n_783, n_784);
  xor g615 (n_785, n_246, n_247);
  xor g616 (n_265, n_785, n_248);
  nand g617 (n_786, n_246, n_247);
  nand g618 (n_787, n_248, n_247);
  nand g619 (n_788, n_246, n_248);
  nand g620 (n_322, n_786, n_787, n_788);
  xor g621 (n_789, n_249, n_250);
  xor g622 (n_270, n_789, n_251);
  nand g623 (n_790, n_249, n_250);
  nand g624 (n_791, n_251, n_250);
  nand g625 (n_792, n_249, n_251);
  nand g626 (n_324, n_790, n_791, n_792);
  xor g627 (n_793, n_252, n_253);
  xor g628 (n_266, n_793, n_254);
  nand g629 (n_794, n_252, n_253);
  nand g630 (n_795, n_254, n_253);
  nand g631 (n_796, n_252, n_254);
  nand g632 (n_323, n_794, n_795, n_796);
  xor g633 (n_797, n_255, n_256);
  xor g634 (n_272, n_797, n_257);
  nand g635 (n_798, n_255, n_256);
  nand g636 (n_799, n_257, n_256);
  nand g637 (n_800, n_255, n_257);
  nand g638 (n_327, n_798, n_799, n_800);
  xor g639 (n_801, n_258, n_259);
  xor g640 (n_271, n_801, n_260);
  nand g641 (n_802, n_258, n_259);
  nand g642 (n_803, n_260, n_259);
  nand g643 (n_804, n_258, n_260);
  nand g644 (n_325, n_802, n_803, n_804);
  xor g645 (n_805, n_261, n_262);
  xor g646 (n_273, n_805, n_263);
  nand g647 (n_806, n_261, n_262);
  nand g648 (n_807, n_263, n_262);
  nand g649 (n_808, n_261, n_263);
  nand g650 (n_333, n_806, n_807, n_808);
  xor g651 (n_809, n_264, n_265);
  xor g652 (n_275, n_809, n_266);
  nand g653 (n_810, n_264, n_265);
  nand g654 (n_811, n_266, n_265);
  nand g655 (n_812, n_264, n_266);
  nand g656 (n_335, n_810, n_811, n_812);
  xor g657 (n_813, n_267, n_268);
  xor g658 (n_277, n_813, n_269);
  nand g659 (n_814, n_267, n_268);
  nand g660 (n_815, n_269, n_268);
  nand g661 (n_816, n_267, n_269);
  nand g662 (n_334, n_814, n_815, n_816);
  xor g663 (n_817, n_270, n_271);
  xor g664 (n_278, n_817, n_272);
  nand g665 (n_818, n_270, n_271);
  nand g666 (n_819, n_272, n_271);
  nand g667 (n_820, n_270, n_272);
  nand g668 (n_337, n_818, n_819, n_820);
  xor g669 (n_821, n_273, n_274);
  xor g670 (n_280, n_821, n_275);
  nand g671 (n_822, n_273, n_274);
  nand g672 (n_823, n_275, n_274);
  nand g673 (n_824, n_273, n_275);
  nand g674 (n_340, n_822, n_823, n_824);
  xor g675 (n_825, n_276, n_277);
  xor g676 (n_98, n_825, n_278);
  nand g677 (n_826, n_276, n_277);
  nand g678 (n_827, n_278, n_277);
  nand g679 (n_828, n_276, n_278);
  nand g680 (n_342, n_826, n_827, n_828);
  xor g681 (n_829, n_279, n_280);
  xor g682 (n_113, n_829, n_281);
  nand g683 (n_830, n_279, n_280);
  nand g684 (n_831, n_281, n_280);
  nand g685 (n_832, n_279, n_281);
  nand g686 (n_97, n_830, n_831, n_832);
  xor g687 (n_833, n_282, n_283);
  xor g688 (n_318, n_833, n_284);
  nand g689 (n_834, n_282, n_283);
  nand g690 (n_835, n_284, n_283);
  nand g691 (n_836, n_282, n_284);
  nand g692 (n_372, n_834, n_835, n_836);
  xor g693 (n_837, n_285, n_286);
  xor g694 (n_315, n_837, n_287);
  nand g695 (n_838, n_285, n_286);
  nand g696 (n_839, n_287, n_286);
  nand g697 (n_840, n_285, n_287);
  nand g698 (n_373, n_838, n_839, n_840);
  xor g699 (n_841, n_288, n_289);
  xor g700 (n_320, n_841, n_290);
  nand g701 (n_842, n_288, n_289);
  nand g702 (n_843, n_290, n_289);
  nand g703 (n_844, n_288, n_290);
  nand g704 (n_374, n_842, n_843, n_844);
  xor g705 (n_845, n_291, n_292);
  xor g706 (n_319, n_845, n_293);
  nand g707 (n_846, n_291, n_292);
  nand g708 (n_847, n_293, n_292);
  nand g709 (n_848, n_291, n_293);
  nand g710 (n_376, n_846, n_847, n_848);
  xor g711 (n_849, n_294, n_295);
  xor g712 (n_316, n_849, n_296);
  nand g713 (n_850, n_294, n_295);
  nand g714 (n_851, n_296, n_295);
  nand g715 (n_852, n_294, n_296);
  nand g716 (n_370, n_850, n_851, n_852);
  xor g717 (n_853, n_297, n_298);
  xor g718 (n_317, n_853, n_299);
  nand g719 (n_854, n_297, n_298);
  nand g720 (n_855, n_299, n_298);
  nand g721 (n_856, n_297, n_299);
  nand g722 (n_377, n_854, n_855, n_856);
  xor g723 (n_857, n_300, n_301);
  xor g724 (n_321, n_857, n_302);
  nand g725 (n_858, n_300, n_301);
  nand g726 (n_859, n_302, n_301);
  nand g727 (n_860, n_300, n_302);
  nand g728 (n_375, n_858, n_859, n_860);
  xor g729 (n_861, n_303, n_304);
  xor g730 (n_314, n_861, n_305);
  nand g731 (n_862, n_303, n_304);
  nand g732 (n_863, n_305, n_304);
  nand g733 (n_864, n_303, n_305);
  nand g734 (n_371, n_862, n_863, n_864);
  xor g735 (n_865, n_306, n_307);
  xor g736 (n_329, n_865, n_308);
  nand g737 (n_866, n_306, n_307);
  nand g738 (n_867, n_308, n_307);
  nand g739 (n_868, n_306, n_308);
  nand g740 (n_385, n_866, n_867, n_868);
  xor g741 (n_869, n_309, n_310);
  xor g742 (n_328, n_869, n_311);
  nand g743 (n_870, n_309, n_310);
  nand g744 (n_871, n_311, n_310);
  nand g745 (n_872, n_309, n_311);
  nand g746 (n_387, n_870, n_871, n_872);
  xor g747 (n_873, n_312, n_313);
  xor g748 (n_326, n_873, n_314);
  nand g749 (n_874, n_312, n_313);
  nand g750 (n_875, n_314, n_313);
  nand g751 (n_876, n_312, n_314);
  nand g752 (n_390, n_874, n_875, n_876);
  xor g753 (n_877, n_315, n_316);
  xor g754 (n_330, n_877, n_317);
  nand g755 (n_878, n_315, n_316);
  nand g756 (n_879, n_317, n_316);
  nand g757 (n_880, n_315, n_317);
  nand g758 (n_391, n_878, n_879, n_880);
  xor g759 (n_881, n_318, n_319);
  xor g760 (n_331, n_881, n_320);
  nand g761 (n_882, n_318, n_319);
  nand g762 (n_883, n_320, n_319);
  nand g763 (n_884, n_318, n_320);
  nand g764 (n_389, n_882, n_883, n_884);
  xor g765 (n_885, n_321, n_322);
  xor g766 (n_332, n_885, n_323);
  nand g767 (n_886, n_321, n_322);
  nand g768 (n_887, n_323, n_322);
  nand g769 (n_888, n_321, n_323);
  nand g770 (n_395, n_886, n_887, n_888);
  xor g771 (n_889, n_324, n_325);
  xor g772 (n_338, n_889, n_326);
  nand g773 (n_890, n_324, n_325);
  nand g774 (n_891, n_326, n_325);
  nand g775 (n_892, n_324, n_326);
  nand g776 (n_397, n_890, n_891, n_892);
  xor g777 (n_893, n_327, n_328);
  xor g778 (n_336, n_893, n_329);
  nand g779 (n_894, n_327, n_328);
  nand g780 (n_895, n_329, n_328);
  nand g781 (n_896, n_327, n_329);
  nand g782 (n_398, n_894, n_895, n_896);
  xor g783 (n_897, n_330, n_331);
  xor g784 (n_339, n_897, n_332);
  nand g785 (n_898, n_330, n_331);
  nand g786 (n_899, n_332, n_331);
  nand g787 (n_900, n_330, n_332);
  nand g788 (n_401, n_898, n_899, n_900);
  xor g789 (n_901, n_333, n_334);
  xor g790 (n_341, n_901, n_335);
  nand g791 (n_902, n_333, n_334);
  nand g792 (n_903, n_335, n_334);
  nand g793 (n_904, n_333, n_335);
  nand g794 (n_403, n_902, n_903, n_904);
  xor g795 (n_905, n_336, n_337);
  xor g796 (n_343, n_905, n_338);
  nand g797 (n_906, n_336, n_337);
  nand g798 (n_907, n_338, n_337);
  nand g799 (n_908, n_336, n_338);
  nand g800 (n_406, n_906, n_907, n_908);
  xor g801 (n_909, n_339, n_340);
  xor g802 (n_344, n_909, n_341);
  nand g803 (n_910, n_339, n_340);
  nand g804 (n_911, n_341, n_340);
  nand g805 (n_912, n_339, n_341);
  nand g806 (n_408, n_910, n_911, n_912);
  xor g807 (n_913, n_342, n_343);
  xor g808 (n_112, n_913, n_344);
  nand g809 (n_914, n_342, n_343);
  nand g810 (n_915, n_344, n_343);
  nand g811 (n_916, n_342, n_344);
  nand g812 (n_96, n_914, n_915, n_916);
  xor g813 (n_369, n_345, n_346);
  and g814 (n_434, n_345, n_346);
  xor g815 (n_917, n_347, n_348);
  xor g816 (n_381, n_917, n_349);
  nand g817 (n_918, n_347, n_348);
  nand g818 (n_919, n_349, n_348);
  nand g819 (n_920, n_347, n_349);
  nand g820 (n_437, n_918, n_919, n_920);
  xor g821 (n_921, n_350, n_351);
  xor g822 (n_384, n_921, n_352);
  nand g823 (n_922, n_350, n_351);
  nand g824 (n_923, n_352, n_351);
  nand g825 (n_924, n_350, n_352);
  nand g826 (n_438, n_922, n_923, n_924);
  xor g827 (n_925, n_353, n_354);
  xor g828 (n_383, n_925, n_355);
  nand g829 (n_926, n_353, n_354);
  nand g830 (n_927, n_355, n_354);
  nand g831 (n_928, n_353, n_355);
  nand g832 (n_439, n_926, n_927, n_928);
  xor g833 (n_929, n_356, n_357);
  xor g834 (n_382, n_929, n_358);
  nand g835 (n_930, n_356, n_357);
  nand g836 (n_931, n_358, n_357);
  nand g837 (n_932, n_356, n_358);
  nand g838 (n_440, n_930, n_931, n_932);
  xor g839 (n_933, n_359, n_360);
  xor g840 (n_379, n_933, n_361);
  nand g841 (n_934, n_359, n_360);
  nand g842 (n_935, n_361, n_360);
  nand g843 (n_936, n_359, n_361);
  nand g844 (n_441, n_934, n_935, n_936);
  xor g845 (n_937, n_362, n_363);
  xor g846 (n_380, n_937, n_364);
  nand g847 (n_938, n_362, n_363);
  nand g848 (n_939, n_364, n_363);
  nand g849 (n_940, n_362, n_364);
  nand g850 (n_436, n_938, n_939, n_940);
  xor g851 (n_941, n_365, n_366);
  xor g852 (n_378, n_941, n_367);
  nand g853 (n_942, n_365, n_366);
  nand g854 (n_943, n_367, n_366);
  nand g855 (n_944, n_365, n_367);
  nand g856 (n_435, n_942, n_943, n_944);
  xor g857 (n_945, n_368, n_369);
  xor g858 (n_386, n_945, n_370);
  nand g859 (n_946, n_368, n_369);
  nand g860 (n_947, n_370, n_369);
  nand g861 (n_948, n_368, n_370);
  nand g862 (n_450, n_946, n_947, n_948);
  xor g863 (n_949, n_371, n_372);
  xor g864 (n_392, n_949, n_373);
  nand g865 (n_950, n_371, n_372);
  nand g866 (n_951, n_373, n_372);
  nand g867 (n_952, n_371, n_373);
  nand g868 (n_451, n_950, n_951, n_952);
  xor g869 (n_953, n_374, n_375);
  xor g870 (n_388, n_953, n_376);
  nand g871 (n_954, n_374, n_375);
  nand g872 (n_955, n_376, n_375);
  nand g873 (n_956, n_374, n_376);
  nand g874 (n_452, n_954, n_955, n_956);
  xor g875 (n_957, n_377, n_378);
  xor g876 (n_393, n_957, n_379);
  nand g877 (n_958, n_377, n_378);
  nand g878 (n_959, n_379, n_378);
  nand g879 (n_960, n_377, n_379);
  nand g880 (n_455, n_958, n_959, n_960);
  xor g881 (n_961, n_380, n_381);
  xor g882 (n_394, n_961, n_382);
  nand g883 (n_962, n_380, n_381);
  nand g884 (n_963, n_382, n_381);
  nand g885 (n_964, n_380, n_382);
  nand g886 (n_454, n_962, n_963, n_964);
  xor g887 (n_965, n_383, n_384);
  xor g888 (n_396, n_965, n_385);
  nand g889 (n_966, n_383, n_384);
  nand g890 (n_967, n_385, n_384);
  nand g891 (n_968, n_383, n_385);
  nand g892 (n_460, n_966, n_967, n_968);
  xor g893 (n_969, n_386, n_387);
  xor g894 (n_399, n_969, n_388);
  nand g895 (n_970, n_386, n_387);
  nand g896 (n_971, n_388, n_387);
  nand g897 (n_972, n_386, n_388);
  nand g898 (n_462, n_970, n_971, n_972);
  xor g899 (n_973, n_389, n_390);
  xor g900 (n_400, n_973, n_391);
  nand g901 (n_974, n_389, n_390);
  nand g902 (n_975, n_391, n_390);
  nand g903 (n_976, n_389, n_391);
  nand g904 (n_461, n_974, n_975, n_976);
  xor g905 (n_977, n_392, n_393);
  xor g906 (n_402, n_977, n_394);
  nand g907 (n_978, n_392, n_393);
  nand g908 (n_979, n_394, n_393);
  nand g909 (n_980, n_392, n_394);
  nand g910 (n_465, n_978, n_979, n_980);
  xor g911 (n_981, n_395, n_396);
  xor g912 (n_404, n_981, n_397);
  nand g913 (n_982, n_395, n_396);
  nand g914 (n_983, n_397, n_396);
  nand g915 (n_984, n_395, n_397);
  nand g916 (n_468, n_982, n_983, n_984);
  xor g917 (n_985, n_398, n_399);
  xor g918 (n_405, n_985, n_400);
  nand g919 (n_986, n_398, n_399);
  nand g920 (n_987, n_400, n_399);
  nand g921 (n_988, n_398, n_400);
  nand g922 (n_469, n_986, n_987, n_988);
  xor g923 (n_989, n_401, n_402);
  xor g924 (n_407, n_989, n_403);
  nand g925 (n_990, n_401, n_402);
  nand g926 (n_991, n_403, n_402);
  nand g927 (n_992, n_401, n_403);
  nand g928 (n_472, n_990, n_991, n_992);
  xor g929 (n_993, n_404, n_405);
  xor g930 (n_409, n_993, n_406);
  nand g931 (n_994, n_404, n_405);
  nand g932 (n_995, n_406, n_405);
  nand g933 (n_996, n_404, n_406);
  nand g934 (n_474, n_994, n_995, n_996);
  xor g935 (n_997, n_407, n_408);
  xor g936 (n_111, n_997, n_409);
  nand g937 (n_998, n_407, n_408);
  nand g938 (n_999, n_409, n_408);
  nand g939 (n_1000, n_407, n_409);
  nand g940 (n_95, n_998, n_999, n_1000);
  xor g941 (n_1001, n_410, n_411);
  xor g942 (n_446, n_1001, n_412);
  nand g943 (n_1002, n_410, n_411);
  nand g944 (n_1003, n_412, n_411);
  nand g945 (n_1004, n_410, n_412);
  nand g946 (n_494, n_1002, n_1003, n_1004);
  xor g947 (n_1005, n_413, n_414);
  xor g948 (n_443, n_1005, n_415);
  nand g949 (n_1006, n_413, n_414);
  nand g950 (n_1007, n_415, n_414);
  nand g951 (n_1008, n_413, n_415);
  nand g952 (n_495, n_1006, n_1007, n_1008);
  xor g953 (n_1009, n_416, n_417);
  xor g954 (n_449, n_1009, n_418);
  nand g955 (n_1010, n_416, n_417);
  nand g956 (n_1011, n_418, n_417);
  nand g957 (n_1012, n_416, n_418);
  nand g958 (n_496, n_1010, n_1011, n_1012);
  xor g959 (n_1013, n_419, n_420);
  xor g960 (n_448, n_1013, n_421);
  nand g961 (n_1014, n_419, n_420);
  nand g962 (n_1015, n_421, n_420);
  nand g963 (n_1016, n_419, n_421);
  nand g964 (n_497, n_1014, n_1015, n_1016);
  xor g965 (n_1017, n_422, n_423);
  xor g966 (n_447, n_1017, n_424);
  nand g967 (n_1018, n_422, n_423);
  nand g968 (n_1019, n_424, n_423);
  nand g969 (n_1020, n_422, n_424);
  nand g970 (n_498, n_1018, n_1019, n_1020);
  xor g971 (n_1021, n_425, n_426);
  xor g972 (n_444, n_1021, n_427);
  nand g973 (n_1022, n_425, n_426);
  nand g974 (n_1023, n_427, n_426);
  nand g975 (n_1024, n_425, n_427);
  nand g976 (n_499, n_1022, n_1023, n_1024);
  xor g977 (n_1025, n_428, n_429);
  xor g978 (n_445, n_1025, n_430);
  nand g979 (n_1026, n_428, n_429);
  nand g980 (n_1027, n_430, n_429);
  nand g981 (n_1028, n_428, n_430);
  nand g982 (n_500, n_1026, n_1027, n_1028);
  xor g983 (n_1029, n_431, n_432);
  xor g984 (n_442, n_1029, n_433);
  nand g985 (n_1030, n_431, n_432);
  nand g986 (n_1031, n_433, n_432);
  nand g987 (n_1032, n_431, n_433);
  nand g988 (n_501, n_1030, n_1031, n_1032);
  xor g989 (n_1033, n_434, n_435);
  xor g990 (n_457, n_1033, n_436);
  nand g991 (n_1034, n_434, n_435);
  nand g992 (n_1035, n_436, n_435);
  nand g993 (n_1036, n_434, n_436);
  nand g994 (n_508, n_1034, n_1035, n_1036);
  xor g995 (n_1037, n_437, n_438);
  xor g996 (n_456, n_1037, n_439);
  nand g997 (n_1038, n_437, n_438);
  nand g998 (n_1039, n_439, n_438);
  nand g999 (n_1040, n_437, n_439);
  nand g1000 (n_509, n_1038, n_1039, n_1040);
  xor g1001 (n_1041, n_440, n_441);
  xor g1002 (n_453, n_1041, n_442);
  nand g1003 (n_1042, n_440, n_441);
  nand g1004 (n_1043, n_442, n_441);
  nand g1005 (n_1044, n_440, n_442);
  nand g1006 (n_513, n_1042, n_1043, n_1044);
  xor g1007 (n_1045, n_443, n_444);
  xor g1008 (n_459, n_1045, n_445);
  nand g1009 (n_1046, n_443, n_444);
  nand g1010 (n_1047, n_445, n_444);
  nand g1011 (n_1048, n_443, n_445);
  nand g1012 (n_515, n_1046, n_1047, n_1048);
  xor g1013 (n_1049, n_446, n_447);
  xor g1014 (n_458, n_1049, n_448);
  nand g1015 (n_1050, n_446, n_447);
  nand g1016 (n_1051, n_448, n_447);
  nand g1017 (n_1052, n_446, n_448);
  nand g1018 (n_512, n_1050, n_1051, n_1052);
  xor g1019 (n_1053, n_449, n_450);
  xor g1020 (n_463, n_1053, n_451);
  nand g1021 (n_1054, n_449, n_450);
  nand g1022 (n_1055, n_451, n_450);
  nand g1023 (n_1056, n_449, n_451);
  nand g1024 (n_517, n_1054, n_1055, n_1056);
  xor g1025 (n_1057, n_452, n_453);
  xor g1026 (n_466, n_1057, n_454);
  nand g1027 (n_1058, n_452, n_453);
  nand g1028 (n_1059, n_454, n_453);
  nand g1029 (n_1060, n_452, n_454);
  nand g1030 (n_520, n_1058, n_1059, n_1060);
  xor g1031 (n_1061, n_455, n_456);
  xor g1032 (n_464, n_1061, n_457);
  nand g1033 (n_1062, n_455, n_456);
  nand g1034 (n_1063, n_457, n_456);
  nand g1035 (n_1064, n_455, n_457);
  nand g1036 (n_519, n_1062, n_1063, n_1064);
  xor g1037 (n_1065, n_458, n_459);
  xor g1038 (n_467, n_1065, n_460);
  nand g1039 (n_1066, n_458, n_459);
  nand g1040 (n_1067, n_460, n_459);
  nand g1041 (n_1068, n_458, n_460);
  nand g1042 (n_524, n_1066, n_1067, n_1068);
  xor g1043 (n_1069, n_461, n_462);
  xor g1044 (n_470, n_1069, n_463);
  nand g1045 (n_1070, n_461, n_462);
  nand g1046 (n_1071, n_463, n_462);
  nand g1047 (n_1072, n_461, n_463);
  nand g1048 (n_525, n_1070, n_1071, n_1072);
  xor g1049 (n_1073, n_464, n_465);
  xor g1050 (n_471, n_1073, n_466);
  nand g1051 (n_1074, n_464, n_465);
  nand g1052 (n_1075, n_466, n_465);
  nand g1053 (n_1076, n_464, n_466);
  nand g1054 (n_526, n_1074, n_1075, n_1076);
  xor g1055 (n_1077, n_467, n_468);
  xor g1056 (n_473, n_1077, n_469);
  nand g1057 (n_1078, n_467, n_468);
  nand g1058 (n_1079, n_469, n_468);
  nand g1059 (n_1080, n_467, n_469);
  nand g1060 (n_529, n_1078, n_1079, n_1080);
  xor g1061 (n_1081, n_470, n_471);
  xor g1062 (n_475, n_1081, n_472);
  nand g1063 (n_1082, n_470, n_471);
  nand g1064 (n_1083, n_472, n_471);
  nand g1065 (n_1084, n_470, n_472);
  nand g1066 (n_531, n_1082, n_1083, n_1084);
  xor g1067 (n_1085, n_473, n_474);
  xor g1068 (n_110, n_1085, n_475);
  nand g1069 (n_1086, n_473, n_474);
  nand g1070 (n_1087, n_475, n_474);
  nand g1071 (n_1088, n_473, n_475);
  nand g1072 (n_94, n_1086, n_1087, n_1088);
  xor g1073 (n_1089, n_476, n_477);
  xor g1074 (n_504, n_1089, n_478);
  nand g1075 (n_1090, n_476, n_477);
  nand g1076 (n_1091, n_478, n_477);
  nand g1077 (n_1092, n_476, n_478);
  nand g1078 (n_550, n_1090, n_1091, n_1092);
  xor g1079 (n_1093, n_479, n_480);
  xor g1080 (n_505, n_1093, n_481);
  nand g1081 (n_1094, n_479, n_480);
  nand g1082 (n_1095, n_481, n_480);
  nand g1083 (n_1096, n_479, n_481);
  nand g1084 (n_551, n_1094, n_1095, n_1096);
  xor g1085 (n_1097, n_482, n_483);
  xor g1086 (n_502, n_1097, n_484);
  nand g1087 (n_1098, n_482, n_483);
  nand g1088 (n_1099, n_484, n_483);
  nand g1089 (n_1100, n_482, n_484);
  nand g1090 (n_546, n_1098, n_1099, n_1100);
  xor g1091 (n_1101, n_485, n_486);
  xor g1092 (n_503, n_1101, n_487);
  nand g1093 (n_1102, n_485, n_486);
  nand g1094 (n_1103, n_487, n_486);
  nand g1095 (n_1104, n_485, n_487);
  nand g1096 (n_547, n_1102, n_1103, n_1104);
  xor g1097 (n_1105, n_488, n_489);
  xor g1098 (n_506, n_1105, n_490);
  nand g1099 (n_1106, n_488, n_489);
  nand g1100 (n_1107, n_490, n_489);
  nand g1101 (n_1108, n_488, n_490);
  nand g1102 (n_548, n_1106, n_1107, n_1108);
  xor g1103 (n_1109, n_491, n_492);
  xor g1104 (n_507, n_1109, n_493);
  nand g1105 (n_1110, n_491, n_492);
  nand g1106 (n_1111, n_493, n_492);
  nand g1107 (n_1112, n_491, n_493);
  nand g1108 (n_549, n_1110, n_1111, n_1112);
  xor g1109 (n_1113, n_494, n_495);
  xor g1110 (n_511, n_1113, n_496);
  nand g1111 (n_1114, n_494, n_495);
  nand g1112 (n_1115, n_496, n_495);
  nand g1113 (n_1116, n_494, n_496);
  nand g1114 (n_555, n_1114, n_1115, n_1116);
  xor g1115 (n_1117, n_497, n_498);
  xor g1116 (n_514, n_1117, n_499);
  nand g1117 (n_1118, n_497, n_498);
  nand g1118 (n_1119, n_499, n_498);
  nand g1119 (n_1120, n_497, n_499);
  nand g1120 (n_556, n_1118, n_1119, n_1120);
  xor g1121 (n_1121, n_500, n_501);
  xor g1122 (n_510, n_1121, n_502);
  nand g1123 (n_1122, n_500, n_501);
  nand g1124 (n_1123, n_502, n_501);
  nand g1125 (n_1124, n_500, n_502);
  nand g1126 (n_560, n_1122, n_1123, n_1124);
  xor g1127 (n_1125, n_503, n_504);
  xor g1128 (n_516, n_1125, n_505);
  nand g1129 (n_1126, n_503, n_504);
  nand g1130 (n_1127, n_505, n_504);
  nand g1131 (n_1128, n_503, n_505);
  nand g1132 (n_558, n_1126, n_1127, n_1128);
  xor g1133 (n_1129, n_506, n_507);
  xor g1134 (n_518, n_1129, n_508);
  nand g1135 (n_1130, n_506, n_507);
  nand g1136 (n_1131, n_508, n_507);
  nand g1137 (n_1132, n_506, n_508);
  nand g1138 (n_562, n_1130, n_1131, n_1132);
  xor g1139 (n_1133, n_509, n_510);
  xor g1140 (n_521, n_1133, n_511);
  nand g1141 (n_1134, n_509, n_510);
  nand g1142 (n_1135, n_511, n_510);
  nand g1143 (n_1136, n_509, n_511);
  nand g1144 (n_565, n_1134, n_1135, n_1136);
  xor g1145 (n_1137, n_512, n_513);
  xor g1146 (n_522, n_1137, n_514);
  nand g1147 (n_1138, n_512, n_513);
  nand g1148 (n_1139, n_514, n_513);
  nand g1149 (n_1140, n_512, n_514);
  nand g1150 (n_566, n_1138, n_1139, n_1140);
  xor g1151 (n_1141, n_515, n_516);
  xor g1152 (n_523, n_1141, n_517);
  nand g1153 (n_1142, n_515, n_516);
  nand g1154 (n_1143, n_517, n_516);
  nand g1155 (n_1144, n_515, n_517);
  nand g1156 (n_568, n_1142, n_1143, n_1144);
  xor g1157 (n_1145, n_518, n_519);
  xor g1158 (n_527, n_1145, n_520);
  nand g1159 (n_1146, n_518, n_519);
  nand g1160 (n_1147, n_520, n_519);
  nand g1161 (n_1148, n_518, n_520);
  nand g1162 (n_569, n_1146, n_1147, n_1148);
  xor g1163 (n_1149, n_521, n_522);
  xor g1164 (n_528, n_1149, n_523);
  nand g1165 (n_1150, n_521, n_522);
  nand g1166 (n_1151, n_523, n_522);
  nand g1167 (n_1152, n_521, n_523);
  nand g1168 (n_572, n_1150, n_1151, n_1152);
  xor g1169 (n_1153, n_524, n_525);
  xor g1170 (n_530, n_1153, n_526);
  nand g1171 (n_1154, n_524, n_525);
  nand g1172 (n_1155, n_526, n_525);
  nand g1173 (n_1156, n_524, n_526);
  nand g1174 (n_573, n_1154, n_1155, n_1156);
  xor g1175 (n_1157, n_527, n_528);
  xor g1176 (n_532, n_1157, n_529);
  nand g1177 (n_1158, n_527, n_528);
  nand g1178 (n_1159, n_529, n_528);
  nand g1179 (n_1160, n_527, n_529);
  nand g1180 (n_576, n_1158, n_1159, n_1160);
  xor g1181 (n_1161, n_530, n_531);
  xor g1182 (n_109, n_1161, n_532);
  nand g1183 (n_1162, n_530, n_531);
  nand g1184 (n_1163, n_532, n_531);
  nand g1185 (n_1164, n_530, n_532);
  nand g1186 (n_93, n_1162, n_1163, n_1164);
  xor g1187 (n_545, n_533, n_534);
  and g1188 (n_584, n_533, n_534);
  xor g1189 (n_1165, n_535, n_536);
  xor g1190 (n_552, n_1165, n_537);
  nand g1191 (n_1166, n_535, n_536);
  nand g1192 (n_1167, n_537, n_536);
  nand g1193 (n_1168, n_535, n_537);
  nand g1194 (n_585, n_1166, n_1167, n_1168);
  xor g1195 (n_1169, n_538, n_539);
  xor g1196 (n_554, n_1169, n_540);
  nand g1197 (n_1170, n_538, n_539);
  nand g1198 (n_1171, n_540, n_539);
  nand g1199 (n_1172, n_538, n_540);
  nand g1200 (n_586, n_1170, n_1171, n_1172);
  xor g1201 (n_1173, n_541, n_542);
  xor g1202 (n_553, n_1173, n_543);
  nand g1203 (n_1174, n_541, n_542);
  nand g1204 (n_1175, n_543, n_542);
  nand g1205 (n_1176, n_541, n_543);
  nand g1206 (n_587, n_1174, n_1175, n_1176);
  xor g1207 (n_1177, n_544, n_545);
  xor g1208 (n_557, n_1177, n_546);
  nand g1209 (n_1178, n_544, n_545);
  nand g1210 (n_1179, n_546, n_545);
  nand g1211 (n_1180, n_544, n_546);
  nand g1212 (n_590, n_1178, n_1179, n_1180);
  xor g1213 (n_1181, n_547, n_548);
  xor g1214 (n_561, n_1181, n_549);
  nand g1215 (n_1182, n_547, n_548);
  nand g1216 (n_1183, n_549, n_548);
  nand g1217 (n_1184, n_547, n_549);
  nand g1218 (n_591, n_1182, n_1183, n_1184);
  xor g1219 (n_1185, n_550, n_551);
  xor g1220 (n_559, n_1185, n_552);
  nand g1221 (n_1186, n_550, n_551);
  nand g1222 (n_1187, n_552, n_551);
  nand g1223 (n_1188, n_550, n_552);
  nand g1224 (n_592, n_1186, n_1187, n_1188);
  xor g1225 (n_1189, n_553, n_554);
  xor g1226 (n_563, n_1189, n_555);
  nand g1227 (n_1190, n_553, n_554);
  nand g1228 (n_1191, n_555, n_554);
  nand g1229 (n_1192, n_553, n_555);
  nand g1230 (n_594, n_1190, n_1191, n_1192);
  xor g1231 (n_1193, n_556, n_557);
  xor g1232 (n_564, n_1193, n_558);
  nand g1233 (n_1194, n_556, n_557);
  nand g1234 (n_1195, n_558, n_557);
  nand g1235 (n_1196, n_556, n_558);
  nand g1236 (n_595, n_1194, n_1195, n_1196);
  xor g1237 (n_1197, n_559, n_560);
  xor g1238 (n_567, n_1197, n_561);
  nand g1239 (n_1198, n_559, n_560);
  nand g1240 (n_1199, n_561, n_560);
  nand g1241 (n_1200, n_559, n_561);
  nand g1242 (n_596, n_1198, n_1199, n_1200);
  xor g1243 (n_1201, n_562, n_563);
  xor g1244 (n_570, n_1201, n_564);
  nand g1245 (n_1202, n_562, n_563);
  nand g1246 (n_1203, n_564, n_563);
  nand g1247 (n_1204, n_562, n_564);
  nand g1248 (n_599, n_1202, n_1203, n_1204);
  xor g1249 (n_1205, n_565, n_566);
  xor g1250 (n_571, n_1205, n_567);
  nand g1251 (n_1206, n_565, n_566);
  nand g1252 (n_1207, n_567, n_566);
  nand g1253 (n_1208, n_565, n_567);
  nand g1254 (n_601, n_1206, n_1207, n_1208);
  xor g1255 (n_1209, n_568, n_569);
  xor g1256 (n_574, n_1209, n_570);
  nand g1257 (n_1210, n_568, n_569);
  nand g1258 (n_1211, n_570, n_569);
  nand g1259 (n_1212, n_568, n_570);
  nand g1260 (n_603, n_1210, n_1211, n_1212);
  xor g1261 (n_1213, n_571, n_572);
  xor g1262 (n_575, n_1213, n_573);
  nand g1263 (n_1214, n_571, n_572);
  nand g1264 (n_1215, n_573, n_572);
  nand g1265 (n_1216, n_571, n_573);
  nand g1266 (n_605, n_1214, n_1215, n_1216);
  xor g1267 (n_1217, n_574, n_575);
  xor g1268 (n_108, n_1217, n_576);
  nand g1269 (n_1218, n_574, n_575);
  nand g1270 (n_1219, n_576, n_575);
  nand g1271 (n_1220, n_574, n_576);
  nand g1272 (n_92, n_1218, n_1219, n_1220);
  xor g1273 (n_583, n_577, n_578);
  and g1274 (n_606, n_577, n_578);
  xor g1275 (n_1221, n_579, n_580);
  xor g1276 (n_588, n_1221, n_581);
  nand g1277 (n_1222, n_579, n_580);
  nand g1278 (n_1223, n_581, n_580);
  nand g1279 (n_1224, n_579, n_581);
  nand g1280 (n_607, n_1222, n_1223, n_1224);
  xor g1281 (n_1225, n_582, n_583);
  xor g1282 (n_589, n_1225, n_584);
  nand g1283 (n_1226, n_582, n_583);
  nand g1284 (n_1227, n_584, n_583);
  nand g1285 (n_1228, n_582, n_584);
  nand g1286 (n_608, n_1226, n_1227, n_1228);
  xor g1287 (n_1229, n_585, n_586);
  xor g1288 (n_593, n_1229, n_587);
  nand g1289 (n_1230, n_585, n_586);
  nand g1290 (n_1231, n_587, n_586);
  nand g1291 (n_1232, n_585, n_587);
  nand g1292 (n_609, n_1230, n_1231, n_1232);
  xor g1293 (n_1233, n_588, n_589);
  xor g1294 (n_597, n_1233, n_590);
  nand g1295 (n_1234, n_588, n_589);
  nand g1296 (n_1235, n_590, n_589);
  nand g1297 (n_1236, n_588, n_590);
  nand g1298 (n_611, n_1234, n_1235, n_1236);
  xor g1299 (n_1237, n_591, n_592);
  xor g1300 (n_598, n_1237, n_593);
  nand g1301 (n_1238, n_591, n_592);
  nand g1302 (n_1239, n_593, n_592);
  nand g1303 (n_1240, n_591, n_593);
  nand g1304 (n_612, n_1238, n_1239, n_1240);
  xor g1305 (n_1241, n_594, n_595);
  xor g1306 (n_600, n_1241, n_596);
  nand g1307 (n_1242, n_594, n_595);
  nand g1308 (n_1243, n_596, n_595);
  nand g1309 (n_1244, n_594, n_596);
  nand g1310 (n_614, n_1242, n_1243, n_1244);
  xor g1311 (n_1245, n_597, n_598);
  xor g1312 (n_602, n_1245, n_599);
  nand g1313 (n_1246, n_597, n_598);
  nand g1314 (n_1247, n_599, n_598);
  nand g1315 (n_1248, n_597, n_599);
  nand g1316 (n_615, n_1246, n_1247, n_1248);
  xor g1317 (n_1249, n_600, n_601);
  xor g1318 (n_604, n_1249, n_602);
  nand g1319 (n_1250, n_600, n_601);
  nand g1320 (n_1251, n_602, n_601);
  nand g1321 (n_1252, n_600, n_602);
  nand g1322 (n_617, n_1250, n_1251, n_1252);
  xor g1323 (n_1253, n_603, n_604);
  xor g1324 (n_107, n_1253, n_605);
  nand g1325 (n_1254, n_603, n_604);
  nand g1326 (n_1255, n_605, n_604);
  nand g1327 (n_1256, n_603, n_605);
  nand g1328 (n_106, n_1254, n_1255, n_1256);
  xor g1329 (n_1257, n_606, n_607);
  xor g1330 (n_610, n_1257, n_608);
  nand g1331 (n_1258, n_606, n_607);
  nand g1332 (n_1259, n_608, n_607);
  nand g1333 (n_1260, n_606, n_608);
  nand g1334 (n_618, n_1258, n_1259, n_1260);
  xor g1335 (n_1261, n_609, n_610);
  xor g1336 (n_613, n_1261, n_611);
  nand g1337 (n_1262, n_609, n_610);
  nand g1338 (n_1263, n_611, n_610);
  nand g1339 (n_1264, n_609, n_611);
  nand g1340 (n_619, n_1262, n_1263, n_1264);
  xor g1341 (n_1265, n_612, n_613);
  xor g1342 (n_616, n_1265, n_614);
  nand g1343 (n_1266, n_612, n_613);
  nand g1344 (n_1267, n_614, n_613);
  nand g1345 (n_1268, n_612, n_614);
  nand g1346 (n_620, n_1266, n_1267, n_1268);
  xor g1347 (n_1269, n_615, n_616);
  xor g1348 (n_91, n_1269, n_617);
  nand g1349 (n_1270, n_615, n_616);
  nand g1350 (n_1271, n_617, n_616);
  nand g1351 (n_1272, n_615, n_617);
  nand g1352 (n_105, n_1270, n_1271, n_1272);
  xor g1353 (n_1273, n_618, n_619);
  xor g1354 (n_90, n_1273, n_620);
  nand g1355 (n_1274, n_618, n_619);
  nand g1356 (n_1275, n_620, n_619);
  nand g1357 (n_1276, n_618, n_620);
  nand g1358 (n_89, n_1274, n_1275, n_1276);
  xor g1359 (n_1363, n_102, n_117);
  nand g1360 (n_1277, n_102, n_117);
  nand g1361 (n_1278, n_102, n_118);
  nand g1362 (n_1279, n_117, n_118);
  nand g1363 (n_1281, n_1277, n_1278, n_1279);
  nor g1364 (n_1280, n_101, n_116);
  nand g1365 (n_1283, n_101, n_116);
  nor g1366 (n_1285, n_100, n_115);
  nand g1367 (n_1288, n_100, n_115);
  nor g1368 (n_1290, n_99, n_114);
  nand g1369 (n_1293, n_99, n_114);
  nor g1370 (n_1295, n_98, n_113);
  nand g1371 (n_1298, n_98, n_113);
  nor g1372 (n_1300, n_97, n_112);
  nand g1373 (n_1303, n_97, n_112);
  nor g1374 (n_1305, n_96, n_111);
  nand g1375 (n_1308, n_96, n_111);
  nor g1376 (n_1310, n_95, n_110);
  nand g1377 (n_1313, n_95, n_110);
  nor g1378 (n_1315, n_94, n_109);
  nand g1379 (n_1318, n_94, n_109);
  nor g1380 (n_1320, n_93, n_108);
  nand g1381 (n_1323, n_93, n_108);
  nor g1382 (n_1325, n_92, n_107);
  nand g1383 (n_1328, n_92, n_107);
  nor g1384 (n_1330, n_91, n_106);
  nand g1385 (n_1333, n_91, n_106);
  nor g1386 (n_1335, n_90, n_105);
  nand g1387 (n_1338, n_90, n_105);
  nand g1394 (n_1286, n_1283, n_1365);
  nand g1397 (n_1291, n_1288, n_1367);
  nand g1400 (n_1296, n_1293, n_1369);
  nand g1403 (n_1301, n_1298, n_1372);
  nand g1406 (n_1306, n_1303, n_1375);
  nand g1409 (n_1311, n_1308, n_1380);
  nand g1412 (n_1316, n_1313, n_1385);
  nand g1415 (n_1321, n_1318, n_1386);
  nand g1418 (n_1326, n_1323, n_1387);
  nand g1421 (n_1331, n_1328, n_1388);
  nand g1424 (n_1336, n_1333, n_1389);
  nand g1427 (n_1341, n_1338, n_1390);
  nand g1429 (n_1344, n_1341, n_89);
  xnor g1433 (out_0[1], n_1281, n_1366);
  xnor g1435 (out_0[2], n_1286, n_1368);
  xnor g1437 (out_0[3], n_1291, n_1370);
  xnor g1439 (out_0[4], n_1296, n_1373);
  xnor g1441 (out_0[5], n_1301, n_1374);
  xnor g1443 (out_0[6], n_1306, n_1376);
  xnor g1445 (out_0[7], n_1311, n_1377);
  xnor g1447 (out_0[8], n_1316, n_1381);
  xnor g1449 (out_0[9], n_1321, n_1382);
  xnor g1451 (out_0[10], n_1326, n_1383);
  xnor g1453 (out_0[11], n_1331, n_1384);
  xnor g1455 (out_0[12], n_1336, n_1379);
  xor g1460 (out_0[0], n_118, n_1363);
  or g1461 (n_1365, n_1280, wc);
  not gc (wc, n_1281);
  or g1462 (n_1366, wc0, n_1280);
  not gc0 (wc0, n_1283);
  or g1463 (n_1367, wc1, n_1285);
  not gc1 (wc1, n_1286);
  or g1464 (n_1368, wc2, n_1285);
  not gc2 (wc2, n_1288);
  or g1465 (n_1369, wc3, n_1290);
  not gc3 (wc3, n_1291);
  or g1466 (n_1370, wc4, n_1290);
  not gc4 (wc4, n_1293);
  or g1468 (n_1372, wc5, n_1295);
  not gc5 (wc5, n_1296);
  or g1469 (n_1373, wc6, n_1295);
  not gc6 (wc6, n_1298);
  or g1470 (n_1374, wc7, n_1300);
  not gc7 (wc7, n_1303);
  or g1471 (n_1375, wc8, n_1300);
  not gc8 (wc8, n_1301);
  or g1472 (n_1376, wc9, n_1305);
  not gc9 (wc9, n_1308);
  or g1473 (n_1377, wc10, n_1310);
  not gc10 (wc10, n_1313);
  or g1475 (n_1379, wc11, n_1335);
  not gc11 (wc11, n_1338);
  or g1476 (n_1380, wc12, n_1305);
  not gc12 (wc12, n_1306);
  or g1477 (n_1381, wc13, n_1315);
  not gc13 (wc13, n_1318);
  or g1478 (n_1382, wc14, n_1320);
  not gc14 (wc14, n_1323);
  or g1479 (n_1383, wc15, n_1325);
  not gc15 (wc15, n_1328);
  or g1480 (n_1384, wc16, n_1330);
  not gc16 (wc16, n_1333);
  or g1481 (n_1385, wc17, n_1310);
  not gc17 (wc17, n_1311);
  or g1482 (n_1386, wc18, n_1315);
  not gc18 (wc18, n_1316);
  or g1483 (n_1387, wc19, n_1320);
  not gc19 (wc19, n_1321);
  or g1484 (n_1388, wc20, n_1325);
  not gc20 (wc20, n_1326);
  or g1485 (n_1389, wc21, n_1330);
  not gc21 (wc21, n_1331);
  or g1486 (n_1390, wc22, n_1335);
  not gc22 (wc22, n_1336);
  xor g1487 (out_0[13], n_89, n_1341);
  not g1488 (out_0[14], n_1344);
endmodule

module csa_tree_add_34_74_group_341_GENERIC(in_0, in_1, in_2, in_3,
     in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, out_0);
  input [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  input [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  output [14:0] out_0;
  wire [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  wire [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  wire [14:0] out_0;
  csa_tree_add_34_74_group_341_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .in_5 (in_5),
       .in_6 (in_6), .in_7 (in_7), .in_8 (in_8), .in_9 (in_9), .in_10
       (in_10), .in_11 (in_11), .out_0 (out_0));
endmodule

module csa_tree_add_35_74_group_343_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( ( ( in_8 * in_9 )  + ( in_10 * in_11 )  )  + ( in_6 * in_7 )  )  + ( in_4 * in_5 )  )  + ( in_2 * in_3 )  )  + ( in_0 * in_1 )  )  ;"
  input [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  input [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  output [14:0] out_0;
  wire [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  wire [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  wire [14:0] out_0;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584;
  wire n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592;
  wire n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672;
  wire n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696;
  wire n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704;
  wire n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760;
  wire n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784;
  wire n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792;
  wire n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800;
  wire n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808;
  wire n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816;
  wire n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832;
  wire n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840;
  wire n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848;
  wire n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856;
  wire n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864;
  wire n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872;
  wire n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880;
  wire n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888;
  wire n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896;
  wire n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904;
  wire n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928;
  wire n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936;
  wire n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944;
  wire n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952;
  wire n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960;
  wire n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968;
  wire n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976;
  wire n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984;
  wire n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992;
  wire n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000;
  wire n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016;
  wire n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048;
  wire n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056;
  wire n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064;
  wire n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088;
  wire n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096;
  wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104;
  wire n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112;
  wire n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120;
  wire n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128;
  wire n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136;
  wire n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144;
  wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152;
  wire n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176;
  wire n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184;
  wire n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264;
  wire n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272;
  wire n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280;
  wire n_1281, n_1283, n_1285, n_1286, n_1288, n_1290, n_1291, n_1293;
  wire n_1295, n_1296, n_1298, n_1300, n_1301, n_1303, n_1305, n_1306;
  wire n_1308, n_1310, n_1311, n_1313, n_1315, n_1316, n_1318, n_1320;
  wire n_1321, n_1323, n_1325, n_1326, n_1328, n_1330, n_1331, n_1333;
  wire n_1335, n_1336, n_1338, n_1341, n_1344, n_1363, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1372, n_1373, n_1374, n_1375;
  wire n_1376, n_1377, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390;
  and g1 (n_119, in_0[0], in_1[0]);
  and g2 (n_124, in_0[1], in_1[0]);
  and g3 (n_142, in_0[2], in_1[0]);
  and g4 (n_173, in_0[3], in_1[0]);
  and g5 (n_223, in_0[4], in_1[0]);
  and g6 (n_282, in_0[5], in_1[0]);
  and g7 (n_345, in_0[6], in_1[0]);
  and g8 (n_410, in_0[7], in_1[0]);
  and g9 (n_125, in_0[0], in_1[1]);
  and g10 (n_143, in_0[1], in_1[1]);
  and g11 (n_174, in_0[2], in_1[1]);
  and g12 (n_224, in_0[3], in_1[1]);
  and g13 (n_283, in_0[4], in_1[1]);
  and g14 (n_346, in_0[5], in_1[1]);
  and g15 (n_411, in_0[6], in_1[1]);
  and g16 (n_476, in_0[7], in_1[1]);
  and g17 (n_151, in_0[0], in_1[2]);
  and g18 (n_189, in_0[1], in_1[2]);
  and g19 (n_239, in_0[2], in_1[2]);
  and g20 (n_298, in_0[3], in_1[2]);
  and g21 (n_361, in_0[4], in_1[2]);
  and g22 (n_426, in_0[5], in_1[2]);
  and g23 (n_477, in_0[6], in_1[2]);
  and g24 (n_533, in_0[7], in_1[2]);
  and g25 (n_175, in_0[0], in_1[3]);
  and g26 (n_225, in_0[1], in_1[3]);
  and g27 (n_284, in_0[2], in_1[3]);
  and g28 (n_347, in_0[3], in_1[3]);
  and g29 (n_412, in_0[4], in_1[3]);
  and g30 (n_487, in_0[5], in_1[3]);
  and g31 (n_534, in_0[6], in_1[3]);
  and g32 (n_577, in_0[7], in_1[3]);
  and g33 (n_122, in_2[0], in_3[0]);
  and g34 (n_133, in_2[1], in_3[0]);
  and g35 (n_144, in_2[2], in_3[0]);
  and g36 (n_182, in_2[3], in_3[0]);
  and g37 (n_232, in_2[4], in_3[0]);
  and g38 (n_291, in_2[5], in_3[0]);
  and g39 (n_354, in_2[6], in_3[0]);
  and g40 (n_419, in_2[7], in_3[0]);
  and g41 (n_126, in_2[0], in_3[1]);
  and g42 (n_104, in_2[1], in_3[1]);
  and g43 (n_190, in_2[2], in_3[1]);
  and g44 (n_240, in_2[3], in_3[1]);
  and g45 (n_299, in_2[4], in_3[1]);
  and g46 (n_362, in_2[5], in_3[1]);
  and g47 (n_427, in_2[6], in_3[1]);
  and g48 (n_478, in_2[7], in_3[1]);
  and g49 (n_152, in_2[0], in_3[2]);
  and g50 (n_194, in_2[1], in_3[2]);
  and g51 (n_244, in_2[2], in_3[2]);
  and g52 (n_303, in_2[3], in_3[2]);
  and g53 (n_366, in_2[4], in_3[2]);
  and g54 (n_431, in_2[5], in_3[2]);
  and g55 (n_484, in_2[6], in_3[2]);
  and g56 (n_541, in_2[7], in_3[2]);
  and g57 (n_176, in_2[0], in_3[3]);
  and g58 (n_226, in_2[1], in_3[3]);
  and g59 (n_285, in_2[2], in_3[3]);
  and g60 (n_348, in_2[3], in_3[3]);
  and g61 (n_413, in_2[4], in_3[3]);
  and g62 (n_488, in_2[5], in_3[3]);
  and g63 (n_535, in_2[6], in_3[3]);
  and g64 (n_578, in_2[7], in_3[3]);
  and g65 (n_118, in_4[0], in_5[0]);
  and g66 (n_132, in_4[1], in_5[0]);
  and g67 (n_157, in_4[2], in_5[0]);
  and g68 (n_179, in_4[3], in_5[0]);
  and g69 (n_229, in_4[4], in_5[0]);
  and g70 (n_288, in_4[5], in_5[0]);
  and g71 (n_351, in_4[6], in_5[0]);
  and g72 (n_416, in_4[7], in_5[0]);
  and g73 (n_134, in_4[0], in_5[1]);
  and g74 (n_145, in_4[1], in_5[1]);
  and g75 (n_183, in_4[2], in_5[1]);
  and g76 (n_233, in_4[3], in_5[1]);
  and g77 (n_292, in_4[4], in_5[1]);
  and g78 (n_355, in_4[5], in_5[1]);
  and g79 (n_420, in_4[6], in_5[1]);
  and g80 (n_491, in_4[7], in_5[1]);
  and g81 (n_148, in_4[0], in_5[2]);
  and g82 (n_186, in_4[1], in_5[2]);
  and g83 (n_236, in_4[2], in_5[2]);
  and g84 (n_295, in_4[3], in_5[2]);
  and g85 (n_358, in_4[4], in_5[2]);
  and g86 (n_423, in_4[5], in_5[2]);
  and g87 (n_479, in_4[6], in_5[2]);
  and g88 (n_538, in_4[7], in_5[2]);
  and g89 (n_191, in_4[0], in_5[3]);
  and g90 (n_241, in_4[1], in_5[3]);
  and g91 (n_300, in_4[2], in_5[3]);
  and g92 (n_363, in_4[3], in_5[3]);
  and g93 (n_428, in_4[4], in_5[3]);
  and g94 (n_482, in_4[5], in_5[3]);
  and g95 (n_542, in_4[6], in_5[3]);
  and g96 (n_581, in_4[7], in_5[3]);
  and g97 (n_123, in_6[0], in_7[0]);
  and g98 (n_135, in_6[1], in_7[0]);
  and g99 (n_149, in_6[2], in_7[0]);
  and g100 (n_193, in_6[3], in_7[0]);
  and g101 (n_243, in_6[4], in_7[0]);
  and g102 (n_302, in_6[5], in_7[0]);
  and g103 (n_365, in_6[6], in_7[0]);
  and g104 (n_430, in_6[7], in_7[0]);
  and g105 (n_128, in_6[0], in_7[1]);
  and g106 (n_150, in_6[1], in_7[1]);
  and g107 (n_195, in_6[2], in_7[1]);
  and g108 (n_245, in_6[3], in_7[1]);
  and g109 (n_304, in_6[4], in_7[1]);
  and g110 (n_367, in_6[5], in_7[1]);
  and g111 (n_432, in_6[6], in_7[1]);
  and g112 (n_485, in_6[7], in_7[1]);
  and g113 (n_153, in_6[0], in_7[2]);
  and g114 (n_196, in_6[1], in_7[2]);
  and g115 (n_246, in_6[2], in_7[2]);
  and g116 (n_305, in_6[3], in_7[2]);
  and g117 (n_368, in_6[4], in_7[2]);
  and g118 (n_433, in_6[5], in_7[2]);
  and g119 (n_486, in_6[6], in_7[2]);
  and g120 (n_544, in_6[7], in_7[2]);
  and g121 (n_177, in_6[0], in_7[3]);
  and g122 (n_227, in_6[1], in_7[3]);
  and g123 (n_286, in_6[2], in_7[3]);
  and g124 (n_349, in_6[3], in_7[3]);
  and g125 (n_414, in_6[4], in_7[3]);
  and g126 (n_489, in_6[5], in_7[3]);
  and g127 (n_536, in_6[6], in_7[3]);
  and g128 (n_579, in_6[7], in_7[3]);
  and g129 (n_121, in_8[0], in_9[0]);
  and g130 (n_131, in_8[1], in_9[0]);
  and g131 (n_156, in_8[2], in_9[0]);
  and g132 (n_178, in_8[3], in_9[0]);
  and g133 (n_228, in_8[4], in_9[0]);
  and g134 (n_287, in_8[5], in_9[0]);
  and g135 (n_350, in_8[6], in_9[0]);
  and g136 (n_415, in_8[7], in_9[0]);
  and g137 (n_130, in_8[0], in_9[1]);
  and g138 (n_155, in_8[1], in_9[1]);
  and g139 (n_180, in_8[2], in_9[1]);
  and g140 (n_230, in_8[3], in_9[1]);
  and g141 (n_289, in_8[4], in_9[1]);
  and g142 (n_352, in_8[5], in_9[1]);
  and g143 (n_417, in_8[6], in_9[1]);
  and g144 (n_490, in_8[7], in_9[1]);
  and g145 (n_154, in_8[0], in_9[2]);
  and g146 (n_181, in_8[1], in_9[2]);
  and g147 (n_231, in_8[2], in_9[2]);
  and g148 (n_290, in_8[3], in_9[2]);
  and g149 (n_353, in_8[4], in_9[2]);
  and g150 (n_418, in_8[5], in_9[2]);
  and g151 (n_492, in_8[6], in_9[2]);
  and g152 (n_537, in_8[7], in_9[2]);
  and g153 (n_184, in_8[0], in_9[3]);
  and g154 (n_234, in_8[1], in_9[3]);
  and g155 (n_293, in_8[2], in_9[3]);
  and g156 (n_356, in_8[3], in_9[3]);
  and g157 (n_421, in_8[4], in_9[3]);
  and g158 (n_493, in_8[5], in_9[3]);
  and g159 (n_539, in_8[6], in_9[3]);
  and g160 (n_580, in_8[7], in_9[3]);
  and g161 (n_120, in_10[0], in_11[0]);
  and g162 (n_129, in_10[1], in_11[0]);
  and g163 (n_146, in_10[2], in_11[0]);
  and g164 (n_185, in_10[3], in_11[0]);
  and g165 (n_235, in_10[4], in_11[0]);
  and g166 (n_294, in_10[5], in_11[0]);
  and g167 (n_357, in_10[6], in_11[0]);
  and g168 (n_422, in_10[7], in_11[0]);
  and g169 (n_127, in_10[0], in_11[1]);
  and g170 (n_147, in_10[1], in_11[1]);
  and g171 (n_187, in_10[2], in_11[1]);
  and g172 (n_237, in_10[3], in_11[1]);
  and g173 (n_296, in_10[4], in_11[1]);
  and g174 (n_359, in_10[5], in_11[1]);
  and g175 (n_424, in_10[6], in_11[1]);
  and g176 (n_480, in_10[7], in_11[1]);
  and g177 (n_103, in_10[0], in_11[2]);
  and g178 (n_188, in_10[1], in_11[2]);
  and g179 (n_238, in_10[2], in_11[2]);
  and g180 (n_297, in_10[3], in_11[2]);
  and g181 (n_360, in_10[4], in_11[2]);
  and g182 (n_425, in_10[5], in_11[2]);
  and g183 (n_481, in_10[6], in_11[2]);
  and g184 (n_540, in_10[7], in_11[2]);
  and g185 (n_192, in_10[0], in_11[3]);
  and g186 (n_242, in_10[1], in_11[3]);
  and g187 (n_301, in_10[2], in_11[3]);
  and g188 (n_364, in_10[3], in_11[3]);
  and g189 (n_429, in_10[4], in_11[3]);
  and g190 (n_483, in_10[5], in_11[3]);
  and g191 (n_543, in_10[6], in_11[3]);
  and g192 (n_582, in_10[7], in_11[3]);
  xor g363 (n_102, n_119, n_120);
  and g364 (n_136, n_119, n_120);
  xor g365 (n_621, n_121, n_122);
  xor g366 (n_117, n_621, n_123);
  nand g367 (n_622, n_121, n_122);
  nand g368 (n_623, n_123, n_122);
  nand g369 (n_624, n_121, n_123);
  nand g370 (n_137, n_622, n_623, n_624);
  xor g371 (n_625, n_124, n_125);
  xor g372 (n_139, n_625, n_126);
  nand g373 (n_626, n_124, n_125);
  nand g374 (n_627, n_126, n_125);
  nand g375 (n_628, n_124, n_126);
  nand g376 (n_161, n_626, n_627, n_628);
  xor g377 (n_629, n_127, n_128);
  xor g378 (n_138, n_629, n_129);
  nand g379 (n_630, n_127, n_128);
  nand g380 (n_631, n_129, n_128);
  nand g381 (n_632, n_127, n_129);
  nand g382 (n_158, n_630, n_631, n_632);
  xor g383 (n_633, n_130, n_131);
  xor g384 (n_141, n_633, n_132);
  nand g385 (n_634, n_130, n_131);
  nand g386 (n_635, n_132, n_131);
  nand g387 (n_636, n_130, n_132);
  nand g388 (n_160, n_634, n_635, n_636);
  xor g389 (n_637, n_133, n_134);
  xor g390 (n_140, n_637, n_135);
  nand g391 (n_638, n_133, n_134);
  nand g392 (n_639, n_135, n_134);
  nand g393 (n_640, n_133, n_135);
  nand g394 (n_159, n_638, n_639, n_640);
  xor g395 (n_641, n_136, n_137);
  xor g396 (n_101, n_641, n_138);
  nand g397 (n_642, n_136, n_137);
  nand g398 (n_643, n_138, n_137);
  nand g399 (n_644, n_136, n_138);
  nand g400 (n_169, n_642, n_643, n_644);
  xor g401 (n_645, n_139, n_140);
  xor g402 (n_116, n_645, n_141);
  nand g403 (n_646, n_139, n_140);
  nand g404 (n_647, n_141, n_140);
  nand g405 (n_648, n_139, n_141);
  nand g406 (n_168, n_646, n_647, n_648);
  xor g407 (n_649, n_142, n_143);
  xor g408 (n_164, n_649, n_144);
  nand g409 (n_650, n_142, n_143);
  nand g410 (n_651, n_144, n_143);
  nand g411 (n_652, n_142, n_144);
  nand g412 (n_202, n_650, n_651, n_652);
  xor g413 (n_653, n_145, n_146);
  xor g414 (n_162, n_653, n_147);
  nand g415 (n_654, n_145, n_146);
  nand g416 (n_655, n_147, n_146);
  nand g417 (n_656, n_145, n_147);
  nand g418 (n_198, n_654, n_655, n_656);
  xor g419 (n_657, n_148, n_103);
  xor g420 (n_163, n_657, n_104);
  nand g421 (n_658, n_148, n_103);
  nand g422 (n_659, n_104, n_103);
  nand g423 (n_660, n_148, n_104);
  nand g424 (n_200, n_658, n_659, n_660);
  xor g425 (n_661, n_149, n_150);
  xor g426 (n_165, n_661, n_151);
  nand g427 (n_662, n_149, n_150);
  nand g428 (n_663, n_151, n_150);
  nand g429 (n_664, n_149, n_151);
  nand g430 (n_203, n_662, n_663, n_664);
  xor g431 (n_665, n_152, n_153);
  xor g432 (n_166, n_665, n_154);
  nand g433 (n_666, n_152, n_153);
  nand g434 (n_667, n_154, n_153);
  nand g435 (n_668, n_152, n_154);
  nand g436 (n_199, n_666, n_667, n_668);
  xor g437 (n_669, n_155, n_156);
  xor g438 (n_167, n_669, n_157);
  nand g439 (n_670, n_155, n_156);
  nand g440 (n_671, n_157, n_156);
  nand g441 (n_672, n_155, n_157);
  nand g442 (n_201, n_670, n_671, n_672);
  xor g443 (n_673, n_158, n_159);
  xor g444 (n_170, n_673, n_160);
  nand g445 (n_674, n_158, n_159);
  nand g446 (n_675, n_160, n_159);
  nand g447 (n_676, n_158, n_160);
  nand g448 (n_211, n_674, n_675, n_676);
  xor g449 (n_677, n_161, n_162);
  xor g450 (n_172, n_677, n_163);
  nand g451 (n_678, n_161, n_162);
  nand g452 (n_679, n_163, n_162);
  nand g453 (n_680, n_161, n_163);
  nand g454 (n_215, n_678, n_679, n_680);
  xor g455 (n_681, n_164, n_165);
  xor g456 (n_171, n_681, n_166);
  nand g457 (n_682, n_164, n_165);
  nand g458 (n_683, n_166, n_165);
  nand g459 (n_684, n_164, n_166);
  nand g460 (n_214, n_682, n_683, n_684);
  xor g461 (n_685, n_167, n_168);
  xor g462 (n_100, n_685, n_169);
  nand g463 (n_686, n_167, n_168);
  nand g464 (n_687, n_169, n_168);
  nand g465 (n_688, n_167, n_169);
  nand g466 (n_220, n_686, n_687, n_688);
  xor g467 (n_689, n_170, n_171);
  xor g468 (n_115, n_689, n_172);
  nand g469 (n_690, n_170, n_171);
  nand g470 (n_691, n_172, n_171);
  nand g471 (n_692, n_170, n_172);
  nand g472 (n_221, n_690, n_691, n_692);
  xor g473 (n_197, n_173, n_174);
  and g474 (n_248, n_173, n_174);
  xor g475 (n_693, n_175, n_176);
  xor g476 (n_206, n_693, n_177);
  nand g477 (n_694, n_175, n_176);
  nand g478 (n_695, n_177, n_176);
  nand g479 (n_696, n_175, n_177);
  nand g480 (n_253, n_694, n_695, n_696);
  xor g481 (n_697, n_178, n_179);
  xor g482 (n_210, n_697, n_180);
  nand g483 (n_698, n_178, n_179);
  nand g484 (n_699, n_180, n_179);
  nand g485 (n_700, n_178, n_180);
  nand g486 (n_254, n_698, n_699, n_700);
  xor g487 (n_701, n_181, n_182);
  xor g488 (n_208, n_701, n_183);
  nand g489 (n_702, n_181, n_182);
  nand g490 (n_703, n_183, n_182);
  nand g491 (n_704, n_181, n_183);
  nand g492 (n_255, n_702, n_703, n_704);
  xor g493 (n_705, n_184, n_185);
  xor g494 (n_205, n_705, n_186);
  nand g495 (n_706, n_184, n_185);
  nand g496 (n_707, n_186, n_185);
  nand g497 (n_708, n_184, n_186);
  nand g498 (n_251, n_706, n_707, n_708);
  xor g499 (n_709, n_187, n_188);
  xor g500 (n_209, n_709, n_189);
  nand g501 (n_710, n_187, n_188);
  nand g502 (n_711, n_189, n_188);
  nand g503 (n_712, n_187, n_189);
  nand g504 (n_250, n_710, n_711, n_712);
  xor g505 (n_713, n_190, n_191);
  xor g506 (n_204, n_713, n_192);
  nand g507 (n_714, n_190, n_191);
  nand g508 (n_715, n_192, n_191);
  nand g509 (n_716, n_190, n_192);
  nand g510 (n_252, n_714, n_715, n_716);
  xor g511 (n_717, n_193, n_194);
  xor g512 (n_207, n_717, n_195);
  nand g513 (n_718, n_193, n_194);
  nand g514 (n_719, n_195, n_194);
  nand g515 (n_720, n_193, n_195);
  nand g516 (n_249, n_718, n_719, n_720);
  xor g517 (n_721, n_196, n_197);
  xor g518 (n_212, n_721, n_198);
  nand g519 (n_722, n_196, n_197);
  nand g520 (n_723, n_198, n_197);
  nand g521 (n_724, n_196, n_198);
  nand g522 (n_263, n_722, n_723, n_724);
  xor g523 (n_725, n_199, n_200);
  xor g524 (n_213, n_725, n_201);
  nand g525 (n_726, n_199, n_200);
  nand g526 (n_727, n_201, n_200);
  nand g527 (n_728, n_199, n_201);
  nand g528 (n_264, n_726, n_727, n_728);
  xor g529 (n_729, n_202, n_203);
  xor g530 (n_216, n_729, n_204);
  nand g531 (n_730, n_202, n_203);
  nand g532 (n_731, n_204, n_203);
  nand g533 (n_732, n_202, n_204);
  nand g534 (n_268, n_730, n_731, n_732);
  xor g535 (n_733, n_205, n_206);
  xor g536 (n_218, n_733, n_207);
  nand g537 (n_734, n_205, n_206);
  nand g538 (n_735, n_207, n_206);
  nand g539 (n_736, n_205, n_207);
  nand g540 (n_267, n_734, n_735, n_736);
  xor g541 (n_737, n_208, n_209);
  xor g542 (n_217, n_737, n_210);
  nand g543 (n_738, n_208, n_209);
  nand g544 (n_739, n_210, n_209);
  nand g545 (n_740, n_208, n_210);
  nand g546 (n_269, n_738, n_739, n_740);
  xor g547 (n_741, n_211, n_212);
  xor g548 (n_219, n_741, n_213);
  nand g549 (n_742, n_211, n_212);
  nand g550 (n_743, n_213, n_212);
  nand g551 (n_744, n_211, n_213);
  nand g552 (n_276, n_742, n_743, n_744);
  xor g553 (n_745, n_214, n_215);
  xor g554 (n_222, n_745, n_216);
  nand g555 (n_746, n_214, n_215);
  nand g556 (n_747, n_216, n_215);
  nand g557 (n_748, n_214, n_216);
  nand g558 (n_274, n_746, n_747, n_748);
  xor g559 (n_749, n_217, n_218);
  xor g560 (n_99, n_749, n_219);
  nand g561 (n_750, n_217, n_218);
  nand g562 (n_751, n_219, n_218);
  nand g563 (n_752, n_217, n_219);
  nand g564 (n_279, n_750, n_751, n_752);
  xor g565 (n_753, n_220, n_221);
  xor g566 (n_114, n_753, n_222);
  nand g567 (n_754, n_220, n_221);
  nand g568 (n_755, n_222, n_221);
  nand g569 (n_756, n_220, n_222);
  nand g570 (n_281, n_754, n_755, n_756);
  xor g571 (n_247, n_223, n_224);
  and g572 (n_306, n_223, n_224);
  xor g573 (n_757, n_225, n_226);
  xor g574 (n_261, n_757, n_227);
  nand g575 (n_758, n_225, n_226);
  nand g576 (n_759, n_227, n_226);
  nand g577 (n_760, n_225, n_227);
  nand g578 (n_309, n_758, n_759, n_760);
  xor g579 (n_761, n_228, n_229);
  xor g580 (n_258, n_761, n_230);
  nand g581 (n_762, n_228, n_229);
  nand g582 (n_763, n_230, n_229);
  nand g583 (n_764, n_228, n_230);
  nand g584 (n_310, n_762, n_763, n_764);
  xor g585 (n_765, n_231, n_232);
  xor g586 (n_260, n_765, n_233);
  nand g587 (n_766, n_231, n_232);
  nand g588 (n_767, n_233, n_232);
  nand g589 (n_768, n_231, n_233);
  nand g590 (n_312, n_766, n_767, n_768);
  xor g591 (n_769, n_234, n_235);
  xor g592 (n_259, n_769, n_236);
  nand g593 (n_770, n_234, n_235);
  nand g594 (n_771, n_236, n_235);
  nand g595 (n_772, n_234, n_236);
  nand g596 (n_308, n_770, n_771, n_772);
  xor g597 (n_773, n_237, n_238);
  xor g598 (n_256, n_773, n_239);
  nand g599 (n_774, n_237, n_238);
  nand g600 (n_775, n_239, n_238);
  nand g601 (n_776, n_237, n_239);
  nand g602 (n_313, n_774, n_775, n_776);
  xor g603 (n_777, n_240, n_241);
  xor g604 (n_262, n_777, n_242);
  nand g605 (n_778, n_240, n_241);
  nand g606 (n_779, n_242, n_241);
  nand g607 (n_780, n_240, n_242);
  nand g608 (n_311, n_778, n_779, n_780);
  xor g609 (n_781, n_243, n_244);
  xor g610 (n_257, n_781, n_245);
  nand g611 (n_782, n_243, n_244);
  nand g612 (n_783, n_245, n_244);
  nand g613 (n_784, n_243, n_245);
  nand g614 (n_307, n_782, n_783, n_784);
  xor g615 (n_785, n_246, n_247);
  xor g616 (n_265, n_785, n_248);
  nand g617 (n_786, n_246, n_247);
  nand g618 (n_787, n_248, n_247);
  nand g619 (n_788, n_246, n_248);
  nand g620 (n_322, n_786, n_787, n_788);
  xor g621 (n_789, n_249, n_250);
  xor g622 (n_270, n_789, n_251);
  nand g623 (n_790, n_249, n_250);
  nand g624 (n_791, n_251, n_250);
  nand g625 (n_792, n_249, n_251);
  nand g626 (n_324, n_790, n_791, n_792);
  xor g627 (n_793, n_252, n_253);
  xor g628 (n_266, n_793, n_254);
  nand g629 (n_794, n_252, n_253);
  nand g630 (n_795, n_254, n_253);
  nand g631 (n_796, n_252, n_254);
  nand g632 (n_323, n_794, n_795, n_796);
  xor g633 (n_797, n_255, n_256);
  xor g634 (n_272, n_797, n_257);
  nand g635 (n_798, n_255, n_256);
  nand g636 (n_799, n_257, n_256);
  nand g637 (n_800, n_255, n_257);
  nand g638 (n_327, n_798, n_799, n_800);
  xor g639 (n_801, n_258, n_259);
  xor g640 (n_271, n_801, n_260);
  nand g641 (n_802, n_258, n_259);
  nand g642 (n_803, n_260, n_259);
  nand g643 (n_804, n_258, n_260);
  nand g644 (n_325, n_802, n_803, n_804);
  xor g645 (n_805, n_261, n_262);
  xor g646 (n_273, n_805, n_263);
  nand g647 (n_806, n_261, n_262);
  nand g648 (n_807, n_263, n_262);
  nand g649 (n_808, n_261, n_263);
  nand g650 (n_333, n_806, n_807, n_808);
  xor g651 (n_809, n_264, n_265);
  xor g652 (n_275, n_809, n_266);
  nand g653 (n_810, n_264, n_265);
  nand g654 (n_811, n_266, n_265);
  nand g655 (n_812, n_264, n_266);
  nand g656 (n_335, n_810, n_811, n_812);
  xor g657 (n_813, n_267, n_268);
  xor g658 (n_277, n_813, n_269);
  nand g659 (n_814, n_267, n_268);
  nand g660 (n_815, n_269, n_268);
  nand g661 (n_816, n_267, n_269);
  nand g662 (n_334, n_814, n_815, n_816);
  xor g663 (n_817, n_270, n_271);
  xor g664 (n_278, n_817, n_272);
  nand g665 (n_818, n_270, n_271);
  nand g666 (n_819, n_272, n_271);
  nand g667 (n_820, n_270, n_272);
  nand g668 (n_337, n_818, n_819, n_820);
  xor g669 (n_821, n_273, n_274);
  xor g670 (n_280, n_821, n_275);
  nand g671 (n_822, n_273, n_274);
  nand g672 (n_823, n_275, n_274);
  nand g673 (n_824, n_273, n_275);
  nand g674 (n_340, n_822, n_823, n_824);
  xor g675 (n_825, n_276, n_277);
  xor g676 (n_98, n_825, n_278);
  nand g677 (n_826, n_276, n_277);
  nand g678 (n_827, n_278, n_277);
  nand g679 (n_828, n_276, n_278);
  nand g680 (n_342, n_826, n_827, n_828);
  xor g681 (n_829, n_279, n_280);
  xor g682 (n_113, n_829, n_281);
  nand g683 (n_830, n_279, n_280);
  nand g684 (n_831, n_281, n_280);
  nand g685 (n_832, n_279, n_281);
  nand g686 (n_97, n_830, n_831, n_832);
  xor g687 (n_833, n_282, n_283);
  xor g688 (n_318, n_833, n_284);
  nand g689 (n_834, n_282, n_283);
  nand g690 (n_835, n_284, n_283);
  nand g691 (n_836, n_282, n_284);
  nand g692 (n_372, n_834, n_835, n_836);
  xor g693 (n_837, n_285, n_286);
  xor g694 (n_315, n_837, n_287);
  nand g695 (n_838, n_285, n_286);
  nand g696 (n_839, n_287, n_286);
  nand g697 (n_840, n_285, n_287);
  nand g698 (n_373, n_838, n_839, n_840);
  xor g699 (n_841, n_288, n_289);
  xor g700 (n_320, n_841, n_290);
  nand g701 (n_842, n_288, n_289);
  nand g702 (n_843, n_290, n_289);
  nand g703 (n_844, n_288, n_290);
  nand g704 (n_374, n_842, n_843, n_844);
  xor g705 (n_845, n_291, n_292);
  xor g706 (n_319, n_845, n_293);
  nand g707 (n_846, n_291, n_292);
  nand g708 (n_847, n_293, n_292);
  nand g709 (n_848, n_291, n_293);
  nand g710 (n_376, n_846, n_847, n_848);
  xor g711 (n_849, n_294, n_295);
  xor g712 (n_316, n_849, n_296);
  nand g713 (n_850, n_294, n_295);
  nand g714 (n_851, n_296, n_295);
  nand g715 (n_852, n_294, n_296);
  nand g716 (n_370, n_850, n_851, n_852);
  xor g717 (n_853, n_297, n_298);
  xor g718 (n_317, n_853, n_299);
  nand g719 (n_854, n_297, n_298);
  nand g720 (n_855, n_299, n_298);
  nand g721 (n_856, n_297, n_299);
  nand g722 (n_377, n_854, n_855, n_856);
  xor g723 (n_857, n_300, n_301);
  xor g724 (n_321, n_857, n_302);
  nand g725 (n_858, n_300, n_301);
  nand g726 (n_859, n_302, n_301);
  nand g727 (n_860, n_300, n_302);
  nand g728 (n_375, n_858, n_859, n_860);
  xor g729 (n_861, n_303, n_304);
  xor g730 (n_314, n_861, n_305);
  nand g731 (n_862, n_303, n_304);
  nand g732 (n_863, n_305, n_304);
  nand g733 (n_864, n_303, n_305);
  nand g734 (n_371, n_862, n_863, n_864);
  xor g735 (n_865, n_306, n_307);
  xor g736 (n_329, n_865, n_308);
  nand g737 (n_866, n_306, n_307);
  nand g738 (n_867, n_308, n_307);
  nand g739 (n_868, n_306, n_308);
  nand g740 (n_385, n_866, n_867, n_868);
  xor g741 (n_869, n_309, n_310);
  xor g742 (n_328, n_869, n_311);
  nand g743 (n_870, n_309, n_310);
  nand g744 (n_871, n_311, n_310);
  nand g745 (n_872, n_309, n_311);
  nand g746 (n_387, n_870, n_871, n_872);
  xor g747 (n_873, n_312, n_313);
  xor g748 (n_326, n_873, n_314);
  nand g749 (n_874, n_312, n_313);
  nand g750 (n_875, n_314, n_313);
  nand g751 (n_876, n_312, n_314);
  nand g752 (n_390, n_874, n_875, n_876);
  xor g753 (n_877, n_315, n_316);
  xor g754 (n_330, n_877, n_317);
  nand g755 (n_878, n_315, n_316);
  nand g756 (n_879, n_317, n_316);
  nand g757 (n_880, n_315, n_317);
  nand g758 (n_391, n_878, n_879, n_880);
  xor g759 (n_881, n_318, n_319);
  xor g760 (n_331, n_881, n_320);
  nand g761 (n_882, n_318, n_319);
  nand g762 (n_883, n_320, n_319);
  nand g763 (n_884, n_318, n_320);
  nand g764 (n_389, n_882, n_883, n_884);
  xor g765 (n_885, n_321, n_322);
  xor g766 (n_332, n_885, n_323);
  nand g767 (n_886, n_321, n_322);
  nand g768 (n_887, n_323, n_322);
  nand g769 (n_888, n_321, n_323);
  nand g770 (n_395, n_886, n_887, n_888);
  xor g771 (n_889, n_324, n_325);
  xor g772 (n_338, n_889, n_326);
  nand g773 (n_890, n_324, n_325);
  nand g774 (n_891, n_326, n_325);
  nand g775 (n_892, n_324, n_326);
  nand g776 (n_397, n_890, n_891, n_892);
  xor g777 (n_893, n_327, n_328);
  xor g778 (n_336, n_893, n_329);
  nand g779 (n_894, n_327, n_328);
  nand g780 (n_895, n_329, n_328);
  nand g781 (n_896, n_327, n_329);
  nand g782 (n_398, n_894, n_895, n_896);
  xor g783 (n_897, n_330, n_331);
  xor g784 (n_339, n_897, n_332);
  nand g785 (n_898, n_330, n_331);
  nand g786 (n_899, n_332, n_331);
  nand g787 (n_900, n_330, n_332);
  nand g788 (n_401, n_898, n_899, n_900);
  xor g789 (n_901, n_333, n_334);
  xor g790 (n_341, n_901, n_335);
  nand g791 (n_902, n_333, n_334);
  nand g792 (n_903, n_335, n_334);
  nand g793 (n_904, n_333, n_335);
  nand g794 (n_403, n_902, n_903, n_904);
  xor g795 (n_905, n_336, n_337);
  xor g796 (n_343, n_905, n_338);
  nand g797 (n_906, n_336, n_337);
  nand g798 (n_907, n_338, n_337);
  nand g799 (n_908, n_336, n_338);
  nand g800 (n_406, n_906, n_907, n_908);
  xor g801 (n_909, n_339, n_340);
  xor g802 (n_344, n_909, n_341);
  nand g803 (n_910, n_339, n_340);
  nand g804 (n_911, n_341, n_340);
  nand g805 (n_912, n_339, n_341);
  nand g806 (n_408, n_910, n_911, n_912);
  xor g807 (n_913, n_342, n_343);
  xor g808 (n_112, n_913, n_344);
  nand g809 (n_914, n_342, n_343);
  nand g810 (n_915, n_344, n_343);
  nand g811 (n_916, n_342, n_344);
  nand g812 (n_96, n_914, n_915, n_916);
  xor g813 (n_369, n_345, n_346);
  and g814 (n_434, n_345, n_346);
  xor g815 (n_917, n_347, n_348);
  xor g816 (n_381, n_917, n_349);
  nand g817 (n_918, n_347, n_348);
  nand g818 (n_919, n_349, n_348);
  nand g819 (n_920, n_347, n_349);
  nand g820 (n_437, n_918, n_919, n_920);
  xor g821 (n_921, n_350, n_351);
  xor g822 (n_384, n_921, n_352);
  nand g823 (n_922, n_350, n_351);
  nand g824 (n_923, n_352, n_351);
  nand g825 (n_924, n_350, n_352);
  nand g826 (n_438, n_922, n_923, n_924);
  xor g827 (n_925, n_353, n_354);
  xor g828 (n_383, n_925, n_355);
  nand g829 (n_926, n_353, n_354);
  nand g830 (n_927, n_355, n_354);
  nand g831 (n_928, n_353, n_355);
  nand g832 (n_439, n_926, n_927, n_928);
  xor g833 (n_929, n_356, n_357);
  xor g834 (n_382, n_929, n_358);
  nand g835 (n_930, n_356, n_357);
  nand g836 (n_931, n_358, n_357);
  nand g837 (n_932, n_356, n_358);
  nand g838 (n_440, n_930, n_931, n_932);
  xor g839 (n_933, n_359, n_360);
  xor g840 (n_379, n_933, n_361);
  nand g841 (n_934, n_359, n_360);
  nand g842 (n_935, n_361, n_360);
  nand g843 (n_936, n_359, n_361);
  nand g844 (n_441, n_934, n_935, n_936);
  xor g845 (n_937, n_362, n_363);
  xor g846 (n_380, n_937, n_364);
  nand g847 (n_938, n_362, n_363);
  nand g848 (n_939, n_364, n_363);
  nand g849 (n_940, n_362, n_364);
  nand g850 (n_436, n_938, n_939, n_940);
  xor g851 (n_941, n_365, n_366);
  xor g852 (n_378, n_941, n_367);
  nand g853 (n_942, n_365, n_366);
  nand g854 (n_943, n_367, n_366);
  nand g855 (n_944, n_365, n_367);
  nand g856 (n_435, n_942, n_943, n_944);
  xor g857 (n_945, n_368, n_369);
  xor g858 (n_386, n_945, n_370);
  nand g859 (n_946, n_368, n_369);
  nand g860 (n_947, n_370, n_369);
  nand g861 (n_948, n_368, n_370);
  nand g862 (n_450, n_946, n_947, n_948);
  xor g863 (n_949, n_371, n_372);
  xor g864 (n_392, n_949, n_373);
  nand g865 (n_950, n_371, n_372);
  nand g866 (n_951, n_373, n_372);
  nand g867 (n_952, n_371, n_373);
  nand g868 (n_451, n_950, n_951, n_952);
  xor g869 (n_953, n_374, n_375);
  xor g870 (n_388, n_953, n_376);
  nand g871 (n_954, n_374, n_375);
  nand g872 (n_955, n_376, n_375);
  nand g873 (n_956, n_374, n_376);
  nand g874 (n_452, n_954, n_955, n_956);
  xor g875 (n_957, n_377, n_378);
  xor g876 (n_393, n_957, n_379);
  nand g877 (n_958, n_377, n_378);
  nand g878 (n_959, n_379, n_378);
  nand g879 (n_960, n_377, n_379);
  nand g880 (n_455, n_958, n_959, n_960);
  xor g881 (n_961, n_380, n_381);
  xor g882 (n_394, n_961, n_382);
  nand g883 (n_962, n_380, n_381);
  nand g884 (n_963, n_382, n_381);
  nand g885 (n_964, n_380, n_382);
  nand g886 (n_454, n_962, n_963, n_964);
  xor g887 (n_965, n_383, n_384);
  xor g888 (n_396, n_965, n_385);
  nand g889 (n_966, n_383, n_384);
  nand g890 (n_967, n_385, n_384);
  nand g891 (n_968, n_383, n_385);
  nand g892 (n_460, n_966, n_967, n_968);
  xor g893 (n_969, n_386, n_387);
  xor g894 (n_399, n_969, n_388);
  nand g895 (n_970, n_386, n_387);
  nand g896 (n_971, n_388, n_387);
  nand g897 (n_972, n_386, n_388);
  nand g898 (n_462, n_970, n_971, n_972);
  xor g899 (n_973, n_389, n_390);
  xor g900 (n_400, n_973, n_391);
  nand g901 (n_974, n_389, n_390);
  nand g902 (n_975, n_391, n_390);
  nand g903 (n_976, n_389, n_391);
  nand g904 (n_461, n_974, n_975, n_976);
  xor g905 (n_977, n_392, n_393);
  xor g906 (n_402, n_977, n_394);
  nand g907 (n_978, n_392, n_393);
  nand g908 (n_979, n_394, n_393);
  nand g909 (n_980, n_392, n_394);
  nand g910 (n_465, n_978, n_979, n_980);
  xor g911 (n_981, n_395, n_396);
  xor g912 (n_404, n_981, n_397);
  nand g913 (n_982, n_395, n_396);
  nand g914 (n_983, n_397, n_396);
  nand g915 (n_984, n_395, n_397);
  nand g916 (n_468, n_982, n_983, n_984);
  xor g917 (n_985, n_398, n_399);
  xor g918 (n_405, n_985, n_400);
  nand g919 (n_986, n_398, n_399);
  nand g920 (n_987, n_400, n_399);
  nand g921 (n_988, n_398, n_400);
  nand g922 (n_469, n_986, n_987, n_988);
  xor g923 (n_989, n_401, n_402);
  xor g924 (n_407, n_989, n_403);
  nand g925 (n_990, n_401, n_402);
  nand g926 (n_991, n_403, n_402);
  nand g927 (n_992, n_401, n_403);
  nand g928 (n_472, n_990, n_991, n_992);
  xor g929 (n_993, n_404, n_405);
  xor g930 (n_409, n_993, n_406);
  nand g931 (n_994, n_404, n_405);
  nand g932 (n_995, n_406, n_405);
  nand g933 (n_996, n_404, n_406);
  nand g934 (n_474, n_994, n_995, n_996);
  xor g935 (n_997, n_407, n_408);
  xor g936 (n_111, n_997, n_409);
  nand g937 (n_998, n_407, n_408);
  nand g938 (n_999, n_409, n_408);
  nand g939 (n_1000, n_407, n_409);
  nand g940 (n_95, n_998, n_999, n_1000);
  xor g941 (n_1001, n_410, n_411);
  xor g942 (n_446, n_1001, n_412);
  nand g943 (n_1002, n_410, n_411);
  nand g944 (n_1003, n_412, n_411);
  nand g945 (n_1004, n_410, n_412);
  nand g946 (n_494, n_1002, n_1003, n_1004);
  xor g947 (n_1005, n_413, n_414);
  xor g948 (n_443, n_1005, n_415);
  nand g949 (n_1006, n_413, n_414);
  nand g950 (n_1007, n_415, n_414);
  nand g951 (n_1008, n_413, n_415);
  nand g952 (n_495, n_1006, n_1007, n_1008);
  xor g953 (n_1009, n_416, n_417);
  xor g954 (n_449, n_1009, n_418);
  nand g955 (n_1010, n_416, n_417);
  nand g956 (n_1011, n_418, n_417);
  nand g957 (n_1012, n_416, n_418);
  nand g958 (n_496, n_1010, n_1011, n_1012);
  xor g959 (n_1013, n_419, n_420);
  xor g960 (n_448, n_1013, n_421);
  nand g961 (n_1014, n_419, n_420);
  nand g962 (n_1015, n_421, n_420);
  nand g963 (n_1016, n_419, n_421);
  nand g964 (n_497, n_1014, n_1015, n_1016);
  xor g965 (n_1017, n_422, n_423);
  xor g966 (n_447, n_1017, n_424);
  nand g967 (n_1018, n_422, n_423);
  nand g968 (n_1019, n_424, n_423);
  nand g969 (n_1020, n_422, n_424);
  nand g970 (n_498, n_1018, n_1019, n_1020);
  xor g971 (n_1021, n_425, n_426);
  xor g972 (n_444, n_1021, n_427);
  nand g973 (n_1022, n_425, n_426);
  nand g974 (n_1023, n_427, n_426);
  nand g975 (n_1024, n_425, n_427);
  nand g976 (n_499, n_1022, n_1023, n_1024);
  xor g977 (n_1025, n_428, n_429);
  xor g978 (n_445, n_1025, n_430);
  nand g979 (n_1026, n_428, n_429);
  nand g980 (n_1027, n_430, n_429);
  nand g981 (n_1028, n_428, n_430);
  nand g982 (n_500, n_1026, n_1027, n_1028);
  xor g983 (n_1029, n_431, n_432);
  xor g984 (n_442, n_1029, n_433);
  nand g985 (n_1030, n_431, n_432);
  nand g986 (n_1031, n_433, n_432);
  nand g987 (n_1032, n_431, n_433);
  nand g988 (n_501, n_1030, n_1031, n_1032);
  xor g989 (n_1033, n_434, n_435);
  xor g990 (n_457, n_1033, n_436);
  nand g991 (n_1034, n_434, n_435);
  nand g992 (n_1035, n_436, n_435);
  nand g993 (n_1036, n_434, n_436);
  nand g994 (n_508, n_1034, n_1035, n_1036);
  xor g995 (n_1037, n_437, n_438);
  xor g996 (n_456, n_1037, n_439);
  nand g997 (n_1038, n_437, n_438);
  nand g998 (n_1039, n_439, n_438);
  nand g999 (n_1040, n_437, n_439);
  nand g1000 (n_509, n_1038, n_1039, n_1040);
  xor g1001 (n_1041, n_440, n_441);
  xor g1002 (n_453, n_1041, n_442);
  nand g1003 (n_1042, n_440, n_441);
  nand g1004 (n_1043, n_442, n_441);
  nand g1005 (n_1044, n_440, n_442);
  nand g1006 (n_513, n_1042, n_1043, n_1044);
  xor g1007 (n_1045, n_443, n_444);
  xor g1008 (n_459, n_1045, n_445);
  nand g1009 (n_1046, n_443, n_444);
  nand g1010 (n_1047, n_445, n_444);
  nand g1011 (n_1048, n_443, n_445);
  nand g1012 (n_515, n_1046, n_1047, n_1048);
  xor g1013 (n_1049, n_446, n_447);
  xor g1014 (n_458, n_1049, n_448);
  nand g1015 (n_1050, n_446, n_447);
  nand g1016 (n_1051, n_448, n_447);
  nand g1017 (n_1052, n_446, n_448);
  nand g1018 (n_512, n_1050, n_1051, n_1052);
  xor g1019 (n_1053, n_449, n_450);
  xor g1020 (n_463, n_1053, n_451);
  nand g1021 (n_1054, n_449, n_450);
  nand g1022 (n_1055, n_451, n_450);
  nand g1023 (n_1056, n_449, n_451);
  nand g1024 (n_517, n_1054, n_1055, n_1056);
  xor g1025 (n_1057, n_452, n_453);
  xor g1026 (n_466, n_1057, n_454);
  nand g1027 (n_1058, n_452, n_453);
  nand g1028 (n_1059, n_454, n_453);
  nand g1029 (n_1060, n_452, n_454);
  nand g1030 (n_520, n_1058, n_1059, n_1060);
  xor g1031 (n_1061, n_455, n_456);
  xor g1032 (n_464, n_1061, n_457);
  nand g1033 (n_1062, n_455, n_456);
  nand g1034 (n_1063, n_457, n_456);
  nand g1035 (n_1064, n_455, n_457);
  nand g1036 (n_519, n_1062, n_1063, n_1064);
  xor g1037 (n_1065, n_458, n_459);
  xor g1038 (n_467, n_1065, n_460);
  nand g1039 (n_1066, n_458, n_459);
  nand g1040 (n_1067, n_460, n_459);
  nand g1041 (n_1068, n_458, n_460);
  nand g1042 (n_524, n_1066, n_1067, n_1068);
  xor g1043 (n_1069, n_461, n_462);
  xor g1044 (n_470, n_1069, n_463);
  nand g1045 (n_1070, n_461, n_462);
  nand g1046 (n_1071, n_463, n_462);
  nand g1047 (n_1072, n_461, n_463);
  nand g1048 (n_525, n_1070, n_1071, n_1072);
  xor g1049 (n_1073, n_464, n_465);
  xor g1050 (n_471, n_1073, n_466);
  nand g1051 (n_1074, n_464, n_465);
  nand g1052 (n_1075, n_466, n_465);
  nand g1053 (n_1076, n_464, n_466);
  nand g1054 (n_526, n_1074, n_1075, n_1076);
  xor g1055 (n_1077, n_467, n_468);
  xor g1056 (n_473, n_1077, n_469);
  nand g1057 (n_1078, n_467, n_468);
  nand g1058 (n_1079, n_469, n_468);
  nand g1059 (n_1080, n_467, n_469);
  nand g1060 (n_529, n_1078, n_1079, n_1080);
  xor g1061 (n_1081, n_470, n_471);
  xor g1062 (n_475, n_1081, n_472);
  nand g1063 (n_1082, n_470, n_471);
  nand g1064 (n_1083, n_472, n_471);
  nand g1065 (n_1084, n_470, n_472);
  nand g1066 (n_531, n_1082, n_1083, n_1084);
  xor g1067 (n_1085, n_473, n_474);
  xor g1068 (n_110, n_1085, n_475);
  nand g1069 (n_1086, n_473, n_474);
  nand g1070 (n_1087, n_475, n_474);
  nand g1071 (n_1088, n_473, n_475);
  nand g1072 (n_94, n_1086, n_1087, n_1088);
  xor g1073 (n_1089, n_476, n_477);
  xor g1074 (n_504, n_1089, n_478);
  nand g1075 (n_1090, n_476, n_477);
  nand g1076 (n_1091, n_478, n_477);
  nand g1077 (n_1092, n_476, n_478);
  nand g1078 (n_550, n_1090, n_1091, n_1092);
  xor g1079 (n_1093, n_479, n_480);
  xor g1080 (n_505, n_1093, n_481);
  nand g1081 (n_1094, n_479, n_480);
  nand g1082 (n_1095, n_481, n_480);
  nand g1083 (n_1096, n_479, n_481);
  nand g1084 (n_551, n_1094, n_1095, n_1096);
  xor g1085 (n_1097, n_482, n_483);
  xor g1086 (n_502, n_1097, n_484);
  nand g1087 (n_1098, n_482, n_483);
  nand g1088 (n_1099, n_484, n_483);
  nand g1089 (n_1100, n_482, n_484);
  nand g1090 (n_546, n_1098, n_1099, n_1100);
  xor g1091 (n_1101, n_485, n_486);
  xor g1092 (n_503, n_1101, n_487);
  nand g1093 (n_1102, n_485, n_486);
  nand g1094 (n_1103, n_487, n_486);
  nand g1095 (n_1104, n_485, n_487);
  nand g1096 (n_547, n_1102, n_1103, n_1104);
  xor g1097 (n_1105, n_488, n_489);
  xor g1098 (n_506, n_1105, n_490);
  nand g1099 (n_1106, n_488, n_489);
  nand g1100 (n_1107, n_490, n_489);
  nand g1101 (n_1108, n_488, n_490);
  nand g1102 (n_548, n_1106, n_1107, n_1108);
  xor g1103 (n_1109, n_491, n_492);
  xor g1104 (n_507, n_1109, n_493);
  nand g1105 (n_1110, n_491, n_492);
  nand g1106 (n_1111, n_493, n_492);
  nand g1107 (n_1112, n_491, n_493);
  nand g1108 (n_549, n_1110, n_1111, n_1112);
  xor g1109 (n_1113, n_494, n_495);
  xor g1110 (n_511, n_1113, n_496);
  nand g1111 (n_1114, n_494, n_495);
  nand g1112 (n_1115, n_496, n_495);
  nand g1113 (n_1116, n_494, n_496);
  nand g1114 (n_555, n_1114, n_1115, n_1116);
  xor g1115 (n_1117, n_497, n_498);
  xor g1116 (n_514, n_1117, n_499);
  nand g1117 (n_1118, n_497, n_498);
  nand g1118 (n_1119, n_499, n_498);
  nand g1119 (n_1120, n_497, n_499);
  nand g1120 (n_556, n_1118, n_1119, n_1120);
  xor g1121 (n_1121, n_500, n_501);
  xor g1122 (n_510, n_1121, n_502);
  nand g1123 (n_1122, n_500, n_501);
  nand g1124 (n_1123, n_502, n_501);
  nand g1125 (n_1124, n_500, n_502);
  nand g1126 (n_560, n_1122, n_1123, n_1124);
  xor g1127 (n_1125, n_503, n_504);
  xor g1128 (n_516, n_1125, n_505);
  nand g1129 (n_1126, n_503, n_504);
  nand g1130 (n_1127, n_505, n_504);
  nand g1131 (n_1128, n_503, n_505);
  nand g1132 (n_558, n_1126, n_1127, n_1128);
  xor g1133 (n_1129, n_506, n_507);
  xor g1134 (n_518, n_1129, n_508);
  nand g1135 (n_1130, n_506, n_507);
  nand g1136 (n_1131, n_508, n_507);
  nand g1137 (n_1132, n_506, n_508);
  nand g1138 (n_562, n_1130, n_1131, n_1132);
  xor g1139 (n_1133, n_509, n_510);
  xor g1140 (n_521, n_1133, n_511);
  nand g1141 (n_1134, n_509, n_510);
  nand g1142 (n_1135, n_511, n_510);
  nand g1143 (n_1136, n_509, n_511);
  nand g1144 (n_565, n_1134, n_1135, n_1136);
  xor g1145 (n_1137, n_512, n_513);
  xor g1146 (n_522, n_1137, n_514);
  nand g1147 (n_1138, n_512, n_513);
  nand g1148 (n_1139, n_514, n_513);
  nand g1149 (n_1140, n_512, n_514);
  nand g1150 (n_566, n_1138, n_1139, n_1140);
  xor g1151 (n_1141, n_515, n_516);
  xor g1152 (n_523, n_1141, n_517);
  nand g1153 (n_1142, n_515, n_516);
  nand g1154 (n_1143, n_517, n_516);
  nand g1155 (n_1144, n_515, n_517);
  nand g1156 (n_568, n_1142, n_1143, n_1144);
  xor g1157 (n_1145, n_518, n_519);
  xor g1158 (n_527, n_1145, n_520);
  nand g1159 (n_1146, n_518, n_519);
  nand g1160 (n_1147, n_520, n_519);
  nand g1161 (n_1148, n_518, n_520);
  nand g1162 (n_569, n_1146, n_1147, n_1148);
  xor g1163 (n_1149, n_521, n_522);
  xor g1164 (n_528, n_1149, n_523);
  nand g1165 (n_1150, n_521, n_522);
  nand g1166 (n_1151, n_523, n_522);
  nand g1167 (n_1152, n_521, n_523);
  nand g1168 (n_572, n_1150, n_1151, n_1152);
  xor g1169 (n_1153, n_524, n_525);
  xor g1170 (n_530, n_1153, n_526);
  nand g1171 (n_1154, n_524, n_525);
  nand g1172 (n_1155, n_526, n_525);
  nand g1173 (n_1156, n_524, n_526);
  nand g1174 (n_573, n_1154, n_1155, n_1156);
  xor g1175 (n_1157, n_527, n_528);
  xor g1176 (n_532, n_1157, n_529);
  nand g1177 (n_1158, n_527, n_528);
  nand g1178 (n_1159, n_529, n_528);
  nand g1179 (n_1160, n_527, n_529);
  nand g1180 (n_576, n_1158, n_1159, n_1160);
  xor g1181 (n_1161, n_530, n_531);
  xor g1182 (n_109, n_1161, n_532);
  nand g1183 (n_1162, n_530, n_531);
  nand g1184 (n_1163, n_532, n_531);
  nand g1185 (n_1164, n_530, n_532);
  nand g1186 (n_93, n_1162, n_1163, n_1164);
  xor g1187 (n_545, n_533, n_534);
  and g1188 (n_584, n_533, n_534);
  xor g1189 (n_1165, n_535, n_536);
  xor g1190 (n_552, n_1165, n_537);
  nand g1191 (n_1166, n_535, n_536);
  nand g1192 (n_1167, n_537, n_536);
  nand g1193 (n_1168, n_535, n_537);
  nand g1194 (n_585, n_1166, n_1167, n_1168);
  xor g1195 (n_1169, n_538, n_539);
  xor g1196 (n_554, n_1169, n_540);
  nand g1197 (n_1170, n_538, n_539);
  nand g1198 (n_1171, n_540, n_539);
  nand g1199 (n_1172, n_538, n_540);
  nand g1200 (n_586, n_1170, n_1171, n_1172);
  xor g1201 (n_1173, n_541, n_542);
  xor g1202 (n_553, n_1173, n_543);
  nand g1203 (n_1174, n_541, n_542);
  nand g1204 (n_1175, n_543, n_542);
  nand g1205 (n_1176, n_541, n_543);
  nand g1206 (n_587, n_1174, n_1175, n_1176);
  xor g1207 (n_1177, n_544, n_545);
  xor g1208 (n_557, n_1177, n_546);
  nand g1209 (n_1178, n_544, n_545);
  nand g1210 (n_1179, n_546, n_545);
  nand g1211 (n_1180, n_544, n_546);
  nand g1212 (n_590, n_1178, n_1179, n_1180);
  xor g1213 (n_1181, n_547, n_548);
  xor g1214 (n_561, n_1181, n_549);
  nand g1215 (n_1182, n_547, n_548);
  nand g1216 (n_1183, n_549, n_548);
  nand g1217 (n_1184, n_547, n_549);
  nand g1218 (n_591, n_1182, n_1183, n_1184);
  xor g1219 (n_1185, n_550, n_551);
  xor g1220 (n_559, n_1185, n_552);
  nand g1221 (n_1186, n_550, n_551);
  nand g1222 (n_1187, n_552, n_551);
  nand g1223 (n_1188, n_550, n_552);
  nand g1224 (n_592, n_1186, n_1187, n_1188);
  xor g1225 (n_1189, n_553, n_554);
  xor g1226 (n_563, n_1189, n_555);
  nand g1227 (n_1190, n_553, n_554);
  nand g1228 (n_1191, n_555, n_554);
  nand g1229 (n_1192, n_553, n_555);
  nand g1230 (n_594, n_1190, n_1191, n_1192);
  xor g1231 (n_1193, n_556, n_557);
  xor g1232 (n_564, n_1193, n_558);
  nand g1233 (n_1194, n_556, n_557);
  nand g1234 (n_1195, n_558, n_557);
  nand g1235 (n_1196, n_556, n_558);
  nand g1236 (n_595, n_1194, n_1195, n_1196);
  xor g1237 (n_1197, n_559, n_560);
  xor g1238 (n_567, n_1197, n_561);
  nand g1239 (n_1198, n_559, n_560);
  nand g1240 (n_1199, n_561, n_560);
  nand g1241 (n_1200, n_559, n_561);
  nand g1242 (n_596, n_1198, n_1199, n_1200);
  xor g1243 (n_1201, n_562, n_563);
  xor g1244 (n_570, n_1201, n_564);
  nand g1245 (n_1202, n_562, n_563);
  nand g1246 (n_1203, n_564, n_563);
  nand g1247 (n_1204, n_562, n_564);
  nand g1248 (n_599, n_1202, n_1203, n_1204);
  xor g1249 (n_1205, n_565, n_566);
  xor g1250 (n_571, n_1205, n_567);
  nand g1251 (n_1206, n_565, n_566);
  nand g1252 (n_1207, n_567, n_566);
  nand g1253 (n_1208, n_565, n_567);
  nand g1254 (n_601, n_1206, n_1207, n_1208);
  xor g1255 (n_1209, n_568, n_569);
  xor g1256 (n_574, n_1209, n_570);
  nand g1257 (n_1210, n_568, n_569);
  nand g1258 (n_1211, n_570, n_569);
  nand g1259 (n_1212, n_568, n_570);
  nand g1260 (n_603, n_1210, n_1211, n_1212);
  xor g1261 (n_1213, n_571, n_572);
  xor g1262 (n_575, n_1213, n_573);
  nand g1263 (n_1214, n_571, n_572);
  nand g1264 (n_1215, n_573, n_572);
  nand g1265 (n_1216, n_571, n_573);
  nand g1266 (n_605, n_1214, n_1215, n_1216);
  xor g1267 (n_1217, n_574, n_575);
  xor g1268 (n_108, n_1217, n_576);
  nand g1269 (n_1218, n_574, n_575);
  nand g1270 (n_1219, n_576, n_575);
  nand g1271 (n_1220, n_574, n_576);
  nand g1272 (n_92, n_1218, n_1219, n_1220);
  xor g1273 (n_583, n_577, n_578);
  and g1274 (n_606, n_577, n_578);
  xor g1275 (n_1221, n_579, n_580);
  xor g1276 (n_588, n_1221, n_581);
  nand g1277 (n_1222, n_579, n_580);
  nand g1278 (n_1223, n_581, n_580);
  nand g1279 (n_1224, n_579, n_581);
  nand g1280 (n_607, n_1222, n_1223, n_1224);
  xor g1281 (n_1225, n_582, n_583);
  xor g1282 (n_589, n_1225, n_584);
  nand g1283 (n_1226, n_582, n_583);
  nand g1284 (n_1227, n_584, n_583);
  nand g1285 (n_1228, n_582, n_584);
  nand g1286 (n_608, n_1226, n_1227, n_1228);
  xor g1287 (n_1229, n_585, n_586);
  xor g1288 (n_593, n_1229, n_587);
  nand g1289 (n_1230, n_585, n_586);
  nand g1290 (n_1231, n_587, n_586);
  nand g1291 (n_1232, n_585, n_587);
  nand g1292 (n_609, n_1230, n_1231, n_1232);
  xor g1293 (n_1233, n_588, n_589);
  xor g1294 (n_597, n_1233, n_590);
  nand g1295 (n_1234, n_588, n_589);
  nand g1296 (n_1235, n_590, n_589);
  nand g1297 (n_1236, n_588, n_590);
  nand g1298 (n_611, n_1234, n_1235, n_1236);
  xor g1299 (n_1237, n_591, n_592);
  xor g1300 (n_598, n_1237, n_593);
  nand g1301 (n_1238, n_591, n_592);
  nand g1302 (n_1239, n_593, n_592);
  nand g1303 (n_1240, n_591, n_593);
  nand g1304 (n_612, n_1238, n_1239, n_1240);
  xor g1305 (n_1241, n_594, n_595);
  xor g1306 (n_600, n_1241, n_596);
  nand g1307 (n_1242, n_594, n_595);
  nand g1308 (n_1243, n_596, n_595);
  nand g1309 (n_1244, n_594, n_596);
  nand g1310 (n_614, n_1242, n_1243, n_1244);
  xor g1311 (n_1245, n_597, n_598);
  xor g1312 (n_602, n_1245, n_599);
  nand g1313 (n_1246, n_597, n_598);
  nand g1314 (n_1247, n_599, n_598);
  nand g1315 (n_1248, n_597, n_599);
  nand g1316 (n_615, n_1246, n_1247, n_1248);
  xor g1317 (n_1249, n_600, n_601);
  xor g1318 (n_604, n_1249, n_602);
  nand g1319 (n_1250, n_600, n_601);
  nand g1320 (n_1251, n_602, n_601);
  nand g1321 (n_1252, n_600, n_602);
  nand g1322 (n_617, n_1250, n_1251, n_1252);
  xor g1323 (n_1253, n_603, n_604);
  xor g1324 (n_107, n_1253, n_605);
  nand g1325 (n_1254, n_603, n_604);
  nand g1326 (n_1255, n_605, n_604);
  nand g1327 (n_1256, n_603, n_605);
  nand g1328 (n_106, n_1254, n_1255, n_1256);
  xor g1329 (n_1257, n_606, n_607);
  xor g1330 (n_610, n_1257, n_608);
  nand g1331 (n_1258, n_606, n_607);
  nand g1332 (n_1259, n_608, n_607);
  nand g1333 (n_1260, n_606, n_608);
  nand g1334 (n_618, n_1258, n_1259, n_1260);
  xor g1335 (n_1261, n_609, n_610);
  xor g1336 (n_613, n_1261, n_611);
  nand g1337 (n_1262, n_609, n_610);
  nand g1338 (n_1263, n_611, n_610);
  nand g1339 (n_1264, n_609, n_611);
  nand g1340 (n_619, n_1262, n_1263, n_1264);
  xor g1341 (n_1265, n_612, n_613);
  xor g1342 (n_616, n_1265, n_614);
  nand g1343 (n_1266, n_612, n_613);
  nand g1344 (n_1267, n_614, n_613);
  nand g1345 (n_1268, n_612, n_614);
  nand g1346 (n_620, n_1266, n_1267, n_1268);
  xor g1347 (n_1269, n_615, n_616);
  xor g1348 (n_91, n_1269, n_617);
  nand g1349 (n_1270, n_615, n_616);
  nand g1350 (n_1271, n_617, n_616);
  nand g1351 (n_1272, n_615, n_617);
  nand g1352 (n_105, n_1270, n_1271, n_1272);
  xor g1353 (n_1273, n_618, n_619);
  xor g1354 (n_90, n_1273, n_620);
  nand g1355 (n_1274, n_618, n_619);
  nand g1356 (n_1275, n_620, n_619);
  nand g1357 (n_1276, n_618, n_620);
  nand g1358 (n_89, n_1274, n_1275, n_1276);
  xor g1359 (n_1363, n_102, n_117);
  nand g1360 (n_1277, n_102, n_117);
  nand g1361 (n_1278, n_102, n_118);
  nand g1362 (n_1279, n_117, n_118);
  nand g1363 (n_1281, n_1277, n_1278, n_1279);
  nor g1364 (n_1280, n_101, n_116);
  nand g1365 (n_1283, n_101, n_116);
  nor g1366 (n_1285, n_100, n_115);
  nand g1367 (n_1288, n_100, n_115);
  nor g1368 (n_1290, n_99, n_114);
  nand g1369 (n_1293, n_99, n_114);
  nor g1370 (n_1295, n_98, n_113);
  nand g1371 (n_1298, n_98, n_113);
  nor g1372 (n_1300, n_97, n_112);
  nand g1373 (n_1303, n_97, n_112);
  nor g1374 (n_1305, n_96, n_111);
  nand g1375 (n_1308, n_96, n_111);
  nor g1376 (n_1310, n_95, n_110);
  nand g1377 (n_1313, n_95, n_110);
  nor g1378 (n_1315, n_94, n_109);
  nand g1379 (n_1318, n_94, n_109);
  nor g1380 (n_1320, n_93, n_108);
  nand g1381 (n_1323, n_93, n_108);
  nor g1382 (n_1325, n_92, n_107);
  nand g1383 (n_1328, n_92, n_107);
  nor g1384 (n_1330, n_91, n_106);
  nand g1385 (n_1333, n_91, n_106);
  nor g1386 (n_1335, n_90, n_105);
  nand g1387 (n_1338, n_90, n_105);
  nand g1394 (n_1286, n_1283, n_1365);
  nand g1397 (n_1291, n_1288, n_1367);
  nand g1400 (n_1296, n_1293, n_1369);
  nand g1403 (n_1301, n_1298, n_1372);
  nand g1406 (n_1306, n_1303, n_1375);
  nand g1409 (n_1311, n_1308, n_1380);
  nand g1412 (n_1316, n_1313, n_1385);
  nand g1415 (n_1321, n_1318, n_1386);
  nand g1418 (n_1326, n_1323, n_1387);
  nand g1421 (n_1331, n_1328, n_1388);
  nand g1424 (n_1336, n_1333, n_1389);
  nand g1427 (n_1341, n_1338, n_1390);
  nand g1429 (n_1344, n_1341, n_89);
  xnor g1433 (out_0[1], n_1281, n_1366);
  xnor g1435 (out_0[2], n_1286, n_1368);
  xnor g1437 (out_0[3], n_1291, n_1370);
  xnor g1439 (out_0[4], n_1296, n_1373);
  xnor g1441 (out_0[5], n_1301, n_1374);
  xnor g1443 (out_0[6], n_1306, n_1376);
  xnor g1445 (out_0[7], n_1311, n_1377);
  xnor g1447 (out_0[8], n_1316, n_1381);
  xnor g1449 (out_0[9], n_1321, n_1382);
  xnor g1451 (out_0[10], n_1326, n_1383);
  xnor g1453 (out_0[11], n_1331, n_1384);
  xnor g1455 (out_0[12], n_1336, n_1379);
  xor g1460 (out_0[0], n_118, n_1363);
  or g1461 (n_1365, n_1280, wc);
  not gc (wc, n_1281);
  or g1462 (n_1366, wc0, n_1280);
  not gc0 (wc0, n_1283);
  or g1463 (n_1367, wc1, n_1285);
  not gc1 (wc1, n_1286);
  or g1464 (n_1368, wc2, n_1285);
  not gc2 (wc2, n_1288);
  or g1465 (n_1369, wc3, n_1290);
  not gc3 (wc3, n_1291);
  or g1466 (n_1370, wc4, n_1290);
  not gc4 (wc4, n_1293);
  or g1468 (n_1372, wc5, n_1295);
  not gc5 (wc5, n_1296);
  or g1469 (n_1373, wc6, n_1295);
  not gc6 (wc6, n_1298);
  or g1470 (n_1374, wc7, n_1300);
  not gc7 (wc7, n_1303);
  or g1471 (n_1375, wc8, n_1300);
  not gc8 (wc8, n_1301);
  or g1472 (n_1376, wc9, n_1305);
  not gc9 (wc9, n_1308);
  or g1473 (n_1377, wc10, n_1310);
  not gc10 (wc10, n_1313);
  or g1475 (n_1379, wc11, n_1335);
  not gc11 (wc11, n_1338);
  or g1476 (n_1380, wc12, n_1305);
  not gc12 (wc12, n_1306);
  or g1477 (n_1381, wc13, n_1315);
  not gc13 (wc13, n_1318);
  or g1478 (n_1382, wc14, n_1320);
  not gc14 (wc14, n_1323);
  or g1479 (n_1383, wc15, n_1325);
  not gc15 (wc15, n_1328);
  or g1480 (n_1384, wc16, n_1330);
  not gc16 (wc16, n_1333);
  or g1481 (n_1385, wc17, n_1310);
  not gc17 (wc17, n_1311);
  or g1482 (n_1386, wc18, n_1315);
  not gc18 (wc18, n_1316);
  or g1483 (n_1387, wc19, n_1320);
  not gc19 (wc19, n_1321);
  or g1484 (n_1388, wc20, n_1325);
  not gc20 (wc20, n_1326);
  or g1485 (n_1389, wc21, n_1330);
  not gc21 (wc21, n_1331);
  or g1486 (n_1390, wc22, n_1335);
  not gc22 (wc22, n_1336);
  xor g1487 (out_0[13], n_89, n_1341);
  not g1488 (out_0[14], n_1344);
endmodule

module csa_tree_add_35_74_group_343_GENERIC(in_0, in_1, in_2, in_3,
     in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, out_0);
  input [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  input [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  output [14:0] out_0;
  wire [7:0] in_0, in_2, in_4, in_6, in_8, in_10;
  wire [3:0] in_1, in_3, in_5, in_7, in_9, in_11;
  wire [14:0] out_0;
  csa_tree_add_35_74_group_343_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .in_5 (in_5),
       .in_6 (in_6), .in_7 (in_7), .in_8 (in_8), .in_9 (in_9), .in_10
       (in_10), .in_11 (in_11), .out_0 (out_0));
endmodule

module csa_tree_distance0_add1034_group_327_GENERIC_REAL(in_0, in_1,
     out_0);
// synthesis_equation "assign out_0 = ( ( in_0 * in_0 )  + ( in_1 * in_1 )  )  ;"
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_358, n_365, n_366, n_367, n_368, n_370;
  wire n_371, n_372, n_373, n_374, n_376, n_377, n_378, n_379;
  wire n_380, n_382, n_383, n_384, n_385, n_386, n_388, n_389;
  wire n_390, n_391, n_392, n_394, n_395, n_396, n_397, n_398;
  wire n_400, n_401, n_402, n_403, n_404, n_406, n_413, n_414;
  wire n_416, n_418, n_423, n_424, n_426, n_428, n_433, n_434;
  wire n_436, n_438, n_451, n_455, n_456, n_458, n_462, n_464;
  wire n_466, n_468, n_470, n_473, n_480, n_482, n_485, n_486;
  wire n_488, n_489, n_491, n_503, n_505, n_508, n_512, n_514;
  wire n_517, n_520, n_523, n_525, n_528, n_535, n_536, n_539;
  wire n_540, n_542, n_543, n_544, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579;
  and g1 (n_48, in_0[0], in_0[1]);
  and g2 (n_70, in_0[0], in_0[2]);
  and g3 (n_74, in_0[1], in_0[2]);
  and g4 (n_75, in_0[0], in_0[3]);
  and g5 (n_78, in_0[1], in_0[3]);
  and g6 (n_86, in_0[2], in_0[3]);
  and g7 (n_79, in_0[0], in_0[4]);
  and g8 (n_90, in_0[1], in_0[4]);
  and g9 (n_98, in_0[2], in_0[4]);
  and g10 (n_109, in_0[3], in_0[4]);
  and g11 (n_87, in_0[0], in_0[5]);
  and g12 (n_99, in_0[1], in_0[5]);
  and g13 (n_67, in_0[2], in_0[5]);
  and g14 (n_124, in_0[3], in_0[5]);
  and g15 (n_141, in_0[4], in_0[5]);
  and g16 (n_50, in_0[0], in_0[6]);
  and g17 (n_110, in_0[1], in_0[6]);
  and g18 (n_125, in_0[2], in_0[6]);
  and g19 (n_145, in_0[3], in_0[6]);
  and g20 (n_157, in_0[4], in_0[6]);
  and g21 (n_170, in_0[5], in_0[6]);
  and g22 (n_113, in_0[0], in_0[7]);
  and g23 (n_128, in_0[1], in_0[7]);
  and g24 (n_142, in_0[2], in_0[7]);
  and g25 (n_158, in_0[3], in_0[7]);
  and g26 (n_171, in_0[4], in_0[7]);
  and g27 (n_179, in_0[5], in_0[7]);
  and g28 (n_185, in_0[6], in_0[7]);
  and g29 (n_69, in_1[0], in_1[1]);
  and g30 (n_71, in_1[0], in_1[2]);
  and g31 (n_73, in_1[1], in_1[2]);
  and g32 (n_72, in_1[0], in_1[3]);
  and g33 (n_81, in_1[1], in_1[3]);
  and g34 (n_89, in_1[2], in_1[3]);
  and g35 (n_80, in_1[0], in_1[4]);
  and g36 (n_91, in_1[1], in_1[4]);
  and g37 (n_100, in_1[2], in_1[4]);
  and g38 (n_66, in_1[3], in_1[4]);
  and g39 (n_88, in_1[0], in_1[5]);
  and g40 (n_49, in_1[1], in_1[5]);
  and g41 (n_111, in_1[2], in_1[5]);
  and g42 (n_126, in_1[3], in_1[5]);
  and g43 (n_144, in_1[4], in_1[5]);
  and g44 (n_51, in_1[0], in_1[6]);
  and g45 (n_112, in_1[1], in_1[6]);
  and g46 (n_127, in_1[2], in_1[6]);
  and g47 (n_146, in_1[3], in_1[6]);
  and g48 (n_160, in_1[4], in_1[6]);
  and g49 (n_169, in_1[5], in_1[6]);
  and g50 (n_114, in_1[0], in_1[7]);
  and g51 (n_129, in_1[1], in_1[7]);
  and g52 (n_143, in_1[2], in_1[7]);
  and g53 (n_159, in_1[3], in_1[7]);
  and g54 (n_172, in_1[4], in_1[7]);
  and g55 (n_180, in_1[5], in_1[7]);
  and g56 (n_186, in_1[6], in_1[7]);
  xor g106 (n_189, in_0[1], in_1[1]);
  xor g107 (n_65, n_189, n_69);
  nand g108 (n_190, in_0[1], in_1[1]);
  nand g109 (n_191, n_69, in_1[1]);
  nand g110 (n_192, in_0[1], n_69);
  nand g111 (n_64, n_190, n_191, n_192);
  xor g112 (n_47, n_70, n_71);
  and g113 (n_77, n_70, n_71);
  xor g114 (n_76, in_0[2], in_1[2]);
  and g115 (n_82, in_0[2], in_1[2]);
  xor g116 (n_193, n_72, n_73);
  xor g117 (n_46, n_193, n_74);
  nand g118 (n_194, n_72, n_73);
  nand g119 (n_195, n_74, n_73);
  nand g120 (n_196, n_72, n_74);
  nand g121 (n_84, n_194, n_195, n_196);
  xor g122 (n_197, n_75, n_76);
  xor g123 (n_63, n_197, n_77);
  nand g124 (n_198, n_75, n_76);
  nand g125 (n_199, n_77, n_76);
  nand g126 (n_200, n_75, n_77);
  nand g127 (n_45, n_198, n_199, n_200);
  xor g128 (n_83, n_78, n_79);
  and g129 (n_93, n_78, n_79);
  xor g130 (n_201, n_80, n_81);
  xor g131 (n_85, n_201, n_82);
  nand g132 (n_202, n_80, n_81);
  nand g133 (n_203, n_82, n_81);
  nand g134 (n_204, n_80, n_82);
  nand g135 (n_95, n_202, n_203, n_204);
  xor g136 (n_205, n_83, n_84);
  xor g137 (n_62, n_205, n_85);
  nand g138 (n_206, n_83, n_84);
  nand g139 (n_207, n_85, n_84);
  nand g140 (n_208, n_83, n_85);
  nand g141 (n_44, n_206, n_207, n_208);
  xor g142 (n_92, in_0[3], in_1[3]);
  and g143 (n_101, in_0[3], in_1[3]);
  xor g144 (n_209, n_86, n_87);
  xor g145 (n_96, n_209, n_88);
  nand g146 (n_210, n_86, n_87);
  nand g147 (n_211, n_88, n_87);
  nand g148 (n_212, n_86, n_88);
  nand g149 (n_103, n_210, n_211, n_212);
  xor g150 (n_213, n_89, n_90);
  xor g151 (n_94, n_213, n_91);
  nand g152 (n_214, n_89, n_90);
  nand g153 (n_215, n_91, n_90);
  nand g154 (n_216, n_89, n_91);
  nand g155 (n_104, n_214, n_215, n_216);
  xor g156 (n_217, n_92, n_93);
  xor g157 (n_97, n_217, n_94);
  nand g158 (n_218, n_92, n_93);
  nand g159 (n_219, n_94, n_93);
  nand g160 (n_220, n_92, n_94);
  nand g161 (n_108, n_218, n_219, n_220);
  xor g162 (n_221, n_95, n_96);
  xor g163 (n_61, n_221, n_97);
  nand g164 (n_222, n_95, n_96);
  nand g165 (n_223, n_97, n_96);
  nand g166 (n_224, n_95, n_97);
  nand g167 (n_43, n_222, n_223, n_224);
  xor g168 (n_102, n_98, n_99);
  and g169 (n_115, n_98, n_99);
  xor g170 (n_225, n_100, n_49);
  xor g171 (n_105, n_225, n_50);
  nand g172 (n_226, n_100, n_49);
  nand g173 (n_227, n_50, n_49);
  nand g174 (n_228, n_100, n_50);
  nand g175 (n_116, n_226, n_227, n_228);
  xor g176 (n_229, n_51, n_101);
  xor g177 (n_106, n_229, n_102);
  nand g178 (n_230, n_51, n_101);
  nand g179 (n_231, n_102, n_101);
  nand g180 (n_232, n_51, n_102);
  nand g181 (n_120, n_230, n_231, n_232);
  xor g182 (n_233, n_103, n_104);
  xor g183 (n_107, n_233, n_105);
  nand g184 (n_234, n_103, n_104);
  nand g185 (n_235, n_105, n_104);
  nand g186 (n_236, n_103, n_105);
  nand g187 (n_121, n_234, n_235, n_236);
  xor g188 (n_237, n_106, n_107);
  xor g189 (n_60, n_237, n_108);
  nand g190 (n_238, n_106, n_107);
  nand g191 (n_239, n_108, n_107);
  nand g192 (n_240, n_106, n_108);
  nand g193 (n_42, n_238, n_239, n_240);
  xor g194 (n_68, in_0[4], in_1[4]);
  and g195 (n_130, in_0[4], in_1[4]);
  xor g196 (n_241, n_109, n_110);
  xor g197 (n_117, n_241, n_111);
  nand g198 (n_242, n_109, n_110);
  nand g199 (n_243, n_111, n_110);
  nand g200 (n_244, n_109, n_111);
  nand g201 (n_133, n_242, n_243, n_244);
  xor g202 (n_245, n_112, n_113);
  xor g203 (n_119, n_245, n_114);
  nand g204 (n_246, n_112, n_113);
  nand g205 (n_247, n_114, n_113);
  nand g206 (n_248, n_112, n_114);
  nand g207 (n_132, n_246, n_247, n_248);
  xor g208 (n_249, n_66, n_67);
  xor g209 (n_118, n_249, n_68);
  nand g210 (n_250, n_66, n_67);
  nand g211 (n_251, n_68, n_67);
  nand g212 (n_252, n_66, n_68);
  nand g213 (n_134, n_250, n_251, n_252);
  xor g214 (n_253, n_115, n_116);
  xor g215 (n_122, n_253, n_117);
  nand g216 (n_254, n_115, n_116);
  nand g217 (n_255, n_117, n_116);
  nand g218 (n_256, n_115, n_117);
  nand g219 (n_138, n_254, n_255, n_256);
  xor g220 (n_257, n_118, n_119);
  xor g221 (n_123, n_257, n_120);
  nand g222 (n_258, n_118, n_119);
  nand g223 (n_259, n_120, n_119);
  nand g224 (n_260, n_118, n_120);
  nand g225 (n_139, n_258, n_259, n_260);
  xor g226 (n_261, n_121, n_122);
  xor g227 (n_59, n_261, n_123);
  nand g228 (n_262, n_121, n_122);
  nand g229 (n_263, n_123, n_122);
  nand g230 (n_264, n_121, n_123);
  nand g231 (n_41, n_262, n_263, n_264);
  xor g232 (n_131, n_124, n_125);
  and g233 (n_147, n_124, n_125);
  xor g234 (n_265, n_126, n_127);
  xor g235 (n_135, n_265, n_128);
  nand g236 (n_266, n_126, n_127);
  nand g237 (n_267, n_128, n_127);
  nand g238 (n_268, n_126, n_128);
  nand g239 (n_148, n_266, n_267, n_268);
  xor g240 (n_269, n_129, n_130);
  xor g241 (n_136, n_269, n_131);
  nand g242 (n_270, n_129, n_130);
  nand g243 (n_271, n_131, n_130);
  nand g244 (n_272, n_129, n_131);
  nand g245 (n_151, n_270, n_271, n_272);
  xor g246 (n_273, n_132, n_133);
  xor g247 (n_137, n_273, n_134);
  nand g248 (n_274, n_132, n_133);
  nand g249 (n_275, n_134, n_133);
  nand g250 (n_276, n_132, n_134);
  nand g251 (n_154, n_274, n_275, n_276);
  xor g252 (n_277, n_135, n_136);
  xor g253 (n_140, n_277, n_137);
  nand g254 (n_278, n_135, n_136);
  nand g255 (n_279, n_137, n_136);
  nand g256 (n_280, n_135, n_137);
  nand g257 (n_156, n_278, n_279, n_280);
  xor g258 (n_281, n_138, n_139);
  xor g259 (n_58, n_281, n_140);
  nand g260 (n_282, n_138, n_139);
  nand g261 (n_283, n_140, n_139);
  nand g262 (n_284, n_138, n_140);
  nand g263 (n_40, n_282, n_283, n_284);
  xor g264 (n_285, in_0[5], in_1[5]);
  xor g265 (n_149, n_285, n_141);
  nand g266 (n_286, in_0[5], in_1[5]);
  nand g267 (n_287, n_141, in_1[5]);
  nand g268 (n_288, in_0[5], n_141);
  nand g269 (n_161, n_286, n_287, n_288);
  xor g270 (n_289, n_142, n_143);
  xor g271 (n_150, n_289, n_144);
  nand g272 (n_290, n_142, n_143);
  nand g273 (n_291, n_144, n_143);
  nand g274 (n_292, n_142, n_144);
  nand g275 (n_162, n_290, n_291, n_292);
  xor g276 (n_293, n_145, n_146);
  xor g277 (n_152, n_293, n_147);
  nand g278 (n_294, n_145, n_146);
  nand g279 (n_295, n_147, n_146);
  nand g280 (n_296, n_145, n_147);
  nand g281 (n_164, n_294, n_295, n_296);
  xor g282 (n_297, n_148, n_149);
  xor g283 (n_153, n_297, n_150);
  nand g284 (n_298, n_148, n_149);
  nand g285 (n_299, n_150, n_149);
  nand g286 (n_300, n_148, n_150);
  nand g287 (n_165, n_298, n_299, n_300);
  xor g288 (n_301, n_151, n_152);
  xor g289 (n_155, n_301, n_153);
  nand g290 (n_302, n_151, n_152);
  nand g291 (n_303, n_153, n_152);
  nand g292 (n_304, n_151, n_153);
  nand g293 (n_168, n_302, n_303, n_304);
  xor g294 (n_305, n_154, n_155);
  xor g295 (n_57, n_305, n_156);
  nand g296 (n_306, n_154, n_155);
  nand g297 (n_307, n_156, n_155);
  nand g298 (n_308, n_154, n_156);
  nand g299 (n_39, n_306, n_307, n_308);
  xor g300 (n_309, n_157, n_158);
  xor g301 (n_163, n_309, n_159);
  nand g302 (n_310, n_157, n_158);
  nand g303 (n_311, n_159, n_158);
  nand g304 (n_312, n_157, n_159);
  nand g305 (n_174, n_310, n_311, n_312);
  xor g306 (n_313, n_160, n_161);
  xor g307 (n_166, n_313, n_162);
  nand g308 (n_314, n_160, n_161);
  nand g309 (n_315, n_162, n_161);
  nand g310 (n_316, n_160, n_162);
  nand g311 (n_176, n_314, n_315, n_316);
  xor g312 (n_317, n_163, n_164);
  xor g313 (n_167, n_317, n_165);
  nand g314 (n_318, n_163, n_164);
  nand g315 (n_319, n_165, n_164);
  nand g316 (n_320, n_163, n_165);
  nand g317 (n_178, n_318, n_319, n_320);
  xor g318 (n_321, n_166, n_167);
  xor g319 (n_56, n_321, n_168);
  nand g320 (n_322, n_166, n_167);
  nand g321 (n_323, n_168, n_167);
  nand g322 (n_324, n_166, n_168);
  nand g323 (n_38, n_322, n_323, n_324);
  xor g324 (n_325, in_0[6], in_1[6]);
  xor g325 (n_173, n_325, n_169);
  nand g326 (n_326, in_0[6], in_1[6]);
  nand g327 (n_327, n_169, in_1[6]);
  nand g328 (n_328, in_0[6], n_169);
  nand g329 (n_182, n_326, n_327, n_328);
  xor g330 (n_329, n_170, n_171);
  xor g331 (n_175, n_329, n_172);
  nand g332 (n_330, n_170, n_171);
  nand g333 (n_331, n_172, n_171);
  nand g334 (n_332, n_170, n_172);
  nand g335 (n_181, n_330, n_331, n_332);
  xor g336 (n_333, n_173, n_174);
  xor g337 (n_177, n_333, n_175);
  nand g338 (n_334, n_173, n_174);
  nand g339 (n_335, n_175, n_174);
  nand g340 (n_336, n_173, n_175);
  nand g341 (n_184, n_334, n_335, n_336);
  xor g342 (n_337, n_176, n_177);
  xor g343 (n_55, n_337, n_178);
  nand g344 (n_338, n_176, n_177);
  nand g345 (n_339, n_178, n_177);
  nand g346 (n_340, n_176, n_178);
  nand g347 (n_54, n_338, n_339, n_340);
  xor g348 (n_341, n_179, n_180);
  xor g349 (n_183, n_341, n_181);
  nand g350 (n_342, n_179, n_180);
  nand g351 (n_343, n_181, n_180);
  nand g352 (n_344, n_179, n_181);
  nand g353 (n_188, n_342, n_343, n_344);
  xor g354 (n_345, n_182, n_183);
  xor g355 (n_37, n_345, n_184);
  nand g356 (n_346, n_182, n_183);
  nand g357 (n_347, n_184, n_183);
  nand g358 (n_348, n_182, n_184);
  nand g359 (n_53, n_346, n_347, n_348);
  xor g360 (n_349, in_0[7], in_1[7]);
  xor g361 (n_187, n_349, n_185);
  nand g362 (n_350, in_0[7], in_1[7]);
  nand g363 (n_351, n_185, in_1[7]);
  nand g364 (n_352, in_0[7], n_185);
  nand g365 (n_35, n_350, n_351, n_352);
  xor g366 (n_353, n_186, n_187);
  xor g367 (n_36, n_353, n_188);
  nand g368 (n_354, n_186, n_187);
  nand g369 (n_355, n_188, n_187);
  nand g370 (n_356, n_186, n_188);
  nand g371 (n_52, n_354, n_355, n_356);
  nand g374 (n_358, in_1[0], in_0[0]);
  nor g379 (n_370, n_48, n_65);
  nand g380 (n_365, n_48, n_65);
  nor g381 (n_366, n_47, n_64);
  nand g382 (n_367, n_47, n_64);
  nor g383 (n_376, n_46, n_63);
  nand g384 (n_371, n_46, n_63);
  nor g385 (n_372, n_45, n_62);
  nand g386 (n_373, n_45, n_62);
  nor g387 (n_382, n_44, n_61);
  nand g388 (n_377, n_44, n_61);
  nor g389 (n_378, n_43, n_60);
  nand g390 (n_379, n_43, n_60);
  nor g391 (n_388, n_42, n_59);
  nand g392 (n_383, n_42, n_59);
  nor g393 (n_384, n_41, n_58);
  nand g394 (n_385, n_41, n_58);
  nor g395 (n_394, n_40, n_57);
  nand g396 (n_389, n_40, n_57);
  nor g397 (n_390, n_39, n_56);
  nand g398 (n_391, n_39, n_56);
  nor g399 (n_400, n_38, n_55);
  nand g400 (n_395, n_38, n_55);
  nor g401 (n_396, n_37, n_54);
  nand g402 (n_397, n_37, n_54);
  nor g403 (n_406, n_36, n_53);
  nand g404 (n_401, n_36, n_53);
  nor g405 (n_402, n_35, n_52);
  nand g406 (n_403, n_35, n_52);
  nor g412 (n_368, n_365, n_366);
  nor g416 (n_374, n_371, n_372);
  nor g419 (n_416, n_376, n_372);
  nor g420 (n_380, n_377, n_378);
  nor g423 (n_418, n_382, n_378);
  nor g424 (n_386, n_383, n_384);
  nor g427 (n_426, n_388, n_384);
  nor g57 (n_392, n_389, n_390);
  nor g60 (n_428, n_394, n_390);
  nor g61 (n_398, n_395, n_396);
  nor g64 (n_436, n_400, n_396);
  nor g65 (n_404, n_401, n_402);
  nor g68 (n_438, n_406, n_402);
  nor g74 (n_414, n_382, n_413);
  nand g83 (n_451, n_416, n_418);
  nor g84 (n_424, n_394, n_423);
  nand g93 (n_458, n_426, n_428);
  nor g94 (n_434, n_406, n_433);
  nand g103 (n_466, n_436, n_438);
  nand g428 (n_503, n_371, n_543);
  nand g430 (n_505, n_413, n_544);
  nand g433 (n_508, n_550, n_551);
  nand g436 (n_470, n_561, n_562);
  nor g437 (n_456, n_400, n_455);
  nor g440 (n_480, n_400, n_458);
  nor g446 (n_464, n_462, n_455);
  nor g449 (n_486, n_458, n_462);
  nor g450 (n_468, n_466, n_455);
  nor g453 (n_489, n_458, n_466);
  nand g456 (n_512, n_383, n_572);
  nand g457 (n_473, n_426, n_470);
  nand g458 (n_514, n_423, n_473);
  nand g461 (n_517, n_566, n_573);
  nand g464 (n_520, n_455, n_574);
  nand g465 (n_482, n_480, n_470);
  nand g466 (n_523, n_576, n_482);
  nand g467 (n_485, n_569, n_470);
  nand g468 (n_525, n_577, n_485);
  nand g469 (n_488, n_486, n_470);
  nand g470 (n_528, n_578, n_488);
  nand g471 (n_491, n_489, n_470);
  nand g472 (out_0[16], n_579, n_491);
  xnor g485 (out_0[5], n_503, n_546);
  xnor g487 (out_0[6], n_505, n_547);
  xnor g490 (out_0[7], n_508, n_552);
  xnor g492 (out_0[8], n_470, n_553);
  xnor g495 (out_0[9], n_512, n_558);
  xnor g497 (out_0[10], n_514, n_559);
  xnor g500 (out_0[11], n_517, n_563);
  xnor g503 (out_0[12], n_520, n_564);
  xnor g506 (out_0[13], n_523, n_565);
  xnor g508 (out_0[14], n_525, n_554);
  xnor g511 (out_0[15], n_528, n_555);
  xor g514 (out_0[0], in_0[0], in_1[0]);
  not g515 (out_0[1], n_358);
  or g516 (n_535, wc, n_370);
  not gc (wc, n_365);
  and g517 (n_536, wc0, n_367);
  not gc0 (wc0, n_368);
  not g519 (out_0[2], n_535);
  or g520 (n_539, wc1, n_366);
  not gc1 (wc1, n_367);
  or g521 (n_540, wc2, n_376);
  not gc2 (wc2, n_371);
  xor g523 (out_0[3], n_365, n_539);
  and g524 (n_413, wc3, n_373);
  not gc3 (wc3, n_374);
  or g525 (n_542, wc4, n_382);
  not gc4 (wc4, n_416);
  or g526 (n_543, n_376, n_536);
  or g527 (n_544, n_536, wc5);
  not gc5 (wc5, n_416);
  xor g528 (out_0[4], n_536, n_540);
  or g529 (n_546, wc6, n_372);
  not gc6 (wc6, n_373);
  or g530 (n_547, wc7, n_382);
  not gc7 (wc7, n_377);
  and g531 (n_548, wc8, n_379);
  not gc8 (wc8, n_380);
  and g532 (n_549, wc9, n_403);
  not gc9 (wc9, n_404);
  and g533 (n_550, wc10, n_377);
  not gc10 (wc10, n_414);
  or g534 (n_551, n_536, n_542);
  or g535 (n_552, wc11, n_378);
  not gc11 (wc11, n_379);
  or g536 (n_553, wc12, n_388);
  not gc12 (wc12, n_383);
  or g537 (n_554, wc13, n_406);
  not gc13 (wc13, n_401);
  or g538 (n_555, wc14, n_402);
  not gc14 (wc14, n_403);
  and g539 (n_423, wc15, n_385);
  not gc15 (wc15, n_386);
  and g540 (n_556, wc16, n_418);
  not gc16 (wc16, n_413);
  or g541 (n_557, wc17, n_394);
  not gc17 (wc17, n_426);
  or g542 (n_558, wc18, n_384);
  not gc18 (wc18, n_385);
  or g543 (n_559, wc19, n_394);
  not gc19 (wc19, n_389);
  and g544 (n_560, wc20, n_391);
  not gc20 (wc20, n_392);
  and g545 (n_433, wc21, n_397);
  not gc21 (wc21, n_398);
  and g546 (n_561, wc22, n_548);
  not gc22 (wc22, n_556);
  or g547 (n_462, wc23, n_406);
  not gc23 (wc23, n_436);
  or g548 (n_562, n_451, n_536);
  or g549 (n_563, wc24, n_390);
  not gc24 (wc24, n_391);
  or g550 (n_564, wc25, n_400);
  not gc25 (wc25, n_395);
  or g551 (n_565, wc26, n_396);
  not gc26 (wc26, n_397);
  and g552 (n_566, wc27, n_389);
  not gc27 (wc27, n_424);
  and g553 (n_567, wc28, n_428);
  not gc28 (wc28, n_423);
  and g554 (n_568, wc29, n_438);
  not gc29 (wc29, n_433);
  and g555 (n_569, wc30, n_436);
  not gc30 (wc30, n_458);
  and g556 (n_455, wc31, n_560);
  not gc31 (wc31, n_567);
  and g557 (n_570, wc32, n_401);
  not gc32 (wc32, n_434);
  and g558 (n_571, wc33, n_549);
  not gc33 (wc33, n_568);
  or g559 (n_572, wc34, n_388);
  not gc34 (wc34, n_470);
  or g560 (n_573, n_557, wc35);
  not gc35 (wc35, n_470);
  or g561 (n_574, wc36, n_458);
  not gc36 (wc36, n_470);
  and g562 (n_575, wc37, n_436);
  not gc37 (wc37, n_455);
  and g563 (n_576, wc38, n_395);
  not gc38 (wc38, n_456);
  and g564 (n_577, wc39, n_433);
  not gc39 (wc39, n_575);
  and g565 (n_578, n_570, wc40);
  not gc40 (wc40, n_464);
  and g566 (n_579, n_571, wc41);
  not gc41 (wc41, n_468);
endmodule

module csa_tree_distance0_add1034_group_327_GENERIC(in_0, in_1, out_0);
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  csa_tree_distance0_add1034_group_327_GENERIC_REAL g1(.in_0 (in_0),
       .in_1 (in_1), .out_0 (out_0));
endmodule

module csa_tree_distance1_add1033_group_329_GENERIC_REAL(in_0, in_1,
     out_0);
// synthesis_equation "assign out_0 = ( ( in_0 * in_0 )  + ( in_1 * in_1 )  )  ;"
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_358, n_365, n_366, n_367, n_368, n_370;
  wire n_371, n_372, n_373, n_374, n_376, n_377, n_378, n_379;
  wire n_380, n_382, n_383, n_384, n_385, n_386, n_388, n_389;
  wire n_390, n_391, n_392, n_394, n_395, n_396, n_397, n_398;
  wire n_400, n_401, n_402, n_403, n_404, n_406, n_413, n_414;
  wire n_416, n_418, n_423, n_424, n_426, n_428, n_433, n_434;
  wire n_436, n_438, n_451, n_455, n_456, n_458, n_462, n_464;
  wire n_466, n_468, n_470, n_473, n_480, n_482, n_485, n_486;
  wire n_488, n_489, n_491, n_503, n_505, n_508, n_512, n_514;
  wire n_517, n_520, n_523, n_525, n_528, n_535, n_536, n_539;
  wire n_540, n_542, n_543, n_544, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579;
  and g1 (n_48, in_0[0], in_0[1]);
  and g2 (n_70, in_0[0], in_0[2]);
  and g3 (n_74, in_0[1], in_0[2]);
  and g4 (n_75, in_0[0], in_0[3]);
  and g5 (n_78, in_0[1], in_0[3]);
  and g6 (n_86, in_0[2], in_0[3]);
  and g7 (n_79, in_0[0], in_0[4]);
  and g8 (n_90, in_0[1], in_0[4]);
  and g9 (n_98, in_0[2], in_0[4]);
  and g10 (n_109, in_0[3], in_0[4]);
  and g11 (n_87, in_0[0], in_0[5]);
  and g12 (n_99, in_0[1], in_0[5]);
  and g13 (n_67, in_0[2], in_0[5]);
  and g14 (n_124, in_0[3], in_0[5]);
  and g15 (n_141, in_0[4], in_0[5]);
  and g16 (n_50, in_0[0], in_0[6]);
  and g17 (n_110, in_0[1], in_0[6]);
  and g18 (n_125, in_0[2], in_0[6]);
  and g19 (n_145, in_0[3], in_0[6]);
  and g20 (n_157, in_0[4], in_0[6]);
  and g21 (n_170, in_0[5], in_0[6]);
  and g22 (n_113, in_0[0], in_0[7]);
  and g23 (n_128, in_0[1], in_0[7]);
  and g24 (n_142, in_0[2], in_0[7]);
  and g25 (n_158, in_0[3], in_0[7]);
  and g26 (n_171, in_0[4], in_0[7]);
  and g27 (n_179, in_0[5], in_0[7]);
  and g28 (n_185, in_0[6], in_0[7]);
  and g29 (n_69, in_1[0], in_1[1]);
  and g30 (n_71, in_1[0], in_1[2]);
  and g31 (n_73, in_1[1], in_1[2]);
  and g32 (n_72, in_1[0], in_1[3]);
  and g33 (n_81, in_1[1], in_1[3]);
  and g34 (n_89, in_1[2], in_1[3]);
  and g35 (n_80, in_1[0], in_1[4]);
  and g36 (n_91, in_1[1], in_1[4]);
  and g37 (n_100, in_1[2], in_1[4]);
  and g38 (n_66, in_1[3], in_1[4]);
  and g39 (n_88, in_1[0], in_1[5]);
  and g40 (n_49, in_1[1], in_1[5]);
  and g41 (n_111, in_1[2], in_1[5]);
  and g42 (n_126, in_1[3], in_1[5]);
  and g43 (n_144, in_1[4], in_1[5]);
  and g44 (n_51, in_1[0], in_1[6]);
  and g45 (n_112, in_1[1], in_1[6]);
  and g46 (n_127, in_1[2], in_1[6]);
  and g47 (n_146, in_1[3], in_1[6]);
  and g48 (n_160, in_1[4], in_1[6]);
  and g49 (n_169, in_1[5], in_1[6]);
  and g50 (n_114, in_1[0], in_1[7]);
  and g51 (n_129, in_1[1], in_1[7]);
  and g52 (n_143, in_1[2], in_1[7]);
  and g53 (n_159, in_1[3], in_1[7]);
  and g54 (n_172, in_1[4], in_1[7]);
  and g55 (n_180, in_1[5], in_1[7]);
  and g56 (n_186, in_1[6], in_1[7]);
  xor g106 (n_189, in_0[1], in_1[1]);
  xor g107 (n_65, n_189, n_69);
  nand g108 (n_190, in_0[1], in_1[1]);
  nand g109 (n_191, n_69, in_1[1]);
  nand g110 (n_192, in_0[1], n_69);
  nand g111 (n_64, n_190, n_191, n_192);
  xor g112 (n_47, n_70, n_71);
  and g113 (n_77, n_70, n_71);
  xor g114 (n_76, in_0[2], in_1[2]);
  and g115 (n_82, in_0[2], in_1[2]);
  xor g116 (n_193, n_72, n_73);
  xor g117 (n_46, n_193, n_74);
  nand g118 (n_194, n_72, n_73);
  nand g119 (n_195, n_74, n_73);
  nand g120 (n_196, n_72, n_74);
  nand g121 (n_84, n_194, n_195, n_196);
  xor g122 (n_197, n_75, n_76);
  xor g123 (n_63, n_197, n_77);
  nand g124 (n_198, n_75, n_76);
  nand g125 (n_199, n_77, n_76);
  nand g126 (n_200, n_75, n_77);
  nand g127 (n_45, n_198, n_199, n_200);
  xor g128 (n_83, n_78, n_79);
  and g129 (n_93, n_78, n_79);
  xor g130 (n_201, n_80, n_81);
  xor g131 (n_85, n_201, n_82);
  nand g132 (n_202, n_80, n_81);
  nand g133 (n_203, n_82, n_81);
  nand g134 (n_204, n_80, n_82);
  nand g135 (n_95, n_202, n_203, n_204);
  xor g136 (n_205, n_83, n_84);
  xor g137 (n_62, n_205, n_85);
  nand g138 (n_206, n_83, n_84);
  nand g139 (n_207, n_85, n_84);
  nand g140 (n_208, n_83, n_85);
  nand g141 (n_44, n_206, n_207, n_208);
  xor g142 (n_92, in_0[3], in_1[3]);
  and g143 (n_101, in_0[3], in_1[3]);
  xor g144 (n_209, n_86, n_87);
  xor g145 (n_96, n_209, n_88);
  nand g146 (n_210, n_86, n_87);
  nand g147 (n_211, n_88, n_87);
  nand g148 (n_212, n_86, n_88);
  nand g149 (n_103, n_210, n_211, n_212);
  xor g150 (n_213, n_89, n_90);
  xor g151 (n_94, n_213, n_91);
  nand g152 (n_214, n_89, n_90);
  nand g153 (n_215, n_91, n_90);
  nand g154 (n_216, n_89, n_91);
  nand g155 (n_104, n_214, n_215, n_216);
  xor g156 (n_217, n_92, n_93);
  xor g157 (n_97, n_217, n_94);
  nand g158 (n_218, n_92, n_93);
  nand g159 (n_219, n_94, n_93);
  nand g160 (n_220, n_92, n_94);
  nand g161 (n_108, n_218, n_219, n_220);
  xor g162 (n_221, n_95, n_96);
  xor g163 (n_61, n_221, n_97);
  nand g164 (n_222, n_95, n_96);
  nand g165 (n_223, n_97, n_96);
  nand g166 (n_224, n_95, n_97);
  nand g167 (n_43, n_222, n_223, n_224);
  xor g168 (n_102, n_98, n_99);
  and g169 (n_115, n_98, n_99);
  xor g170 (n_225, n_100, n_49);
  xor g171 (n_105, n_225, n_50);
  nand g172 (n_226, n_100, n_49);
  nand g173 (n_227, n_50, n_49);
  nand g174 (n_228, n_100, n_50);
  nand g175 (n_116, n_226, n_227, n_228);
  xor g176 (n_229, n_51, n_101);
  xor g177 (n_106, n_229, n_102);
  nand g178 (n_230, n_51, n_101);
  nand g179 (n_231, n_102, n_101);
  nand g180 (n_232, n_51, n_102);
  nand g181 (n_120, n_230, n_231, n_232);
  xor g182 (n_233, n_103, n_104);
  xor g183 (n_107, n_233, n_105);
  nand g184 (n_234, n_103, n_104);
  nand g185 (n_235, n_105, n_104);
  nand g186 (n_236, n_103, n_105);
  nand g187 (n_121, n_234, n_235, n_236);
  xor g188 (n_237, n_106, n_107);
  xor g189 (n_60, n_237, n_108);
  nand g190 (n_238, n_106, n_107);
  nand g191 (n_239, n_108, n_107);
  nand g192 (n_240, n_106, n_108);
  nand g193 (n_42, n_238, n_239, n_240);
  xor g194 (n_68, in_0[4], in_1[4]);
  and g195 (n_130, in_0[4], in_1[4]);
  xor g196 (n_241, n_109, n_110);
  xor g197 (n_117, n_241, n_111);
  nand g198 (n_242, n_109, n_110);
  nand g199 (n_243, n_111, n_110);
  nand g200 (n_244, n_109, n_111);
  nand g201 (n_133, n_242, n_243, n_244);
  xor g202 (n_245, n_112, n_113);
  xor g203 (n_119, n_245, n_114);
  nand g204 (n_246, n_112, n_113);
  nand g205 (n_247, n_114, n_113);
  nand g206 (n_248, n_112, n_114);
  nand g207 (n_132, n_246, n_247, n_248);
  xor g208 (n_249, n_66, n_67);
  xor g209 (n_118, n_249, n_68);
  nand g210 (n_250, n_66, n_67);
  nand g211 (n_251, n_68, n_67);
  nand g212 (n_252, n_66, n_68);
  nand g213 (n_134, n_250, n_251, n_252);
  xor g214 (n_253, n_115, n_116);
  xor g215 (n_122, n_253, n_117);
  nand g216 (n_254, n_115, n_116);
  nand g217 (n_255, n_117, n_116);
  nand g218 (n_256, n_115, n_117);
  nand g219 (n_138, n_254, n_255, n_256);
  xor g220 (n_257, n_118, n_119);
  xor g221 (n_123, n_257, n_120);
  nand g222 (n_258, n_118, n_119);
  nand g223 (n_259, n_120, n_119);
  nand g224 (n_260, n_118, n_120);
  nand g225 (n_139, n_258, n_259, n_260);
  xor g226 (n_261, n_121, n_122);
  xor g227 (n_59, n_261, n_123);
  nand g228 (n_262, n_121, n_122);
  nand g229 (n_263, n_123, n_122);
  nand g230 (n_264, n_121, n_123);
  nand g231 (n_41, n_262, n_263, n_264);
  xor g232 (n_131, n_124, n_125);
  and g233 (n_147, n_124, n_125);
  xor g234 (n_265, n_126, n_127);
  xor g235 (n_135, n_265, n_128);
  nand g236 (n_266, n_126, n_127);
  nand g237 (n_267, n_128, n_127);
  nand g238 (n_268, n_126, n_128);
  nand g239 (n_148, n_266, n_267, n_268);
  xor g240 (n_269, n_129, n_130);
  xor g241 (n_136, n_269, n_131);
  nand g242 (n_270, n_129, n_130);
  nand g243 (n_271, n_131, n_130);
  nand g244 (n_272, n_129, n_131);
  nand g245 (n_151, n_270, n_271, n_272);
  xor g246 (n_273, n_132, n_133);
  xor g247 (n_137, n_273, n_134);
  nand g248 (n_274, n_132, n_133);
  nand g249 (n_275, n_134, n_133);
  nand g250 (n_276, n_132, n_134);
  nand g251 (n_154, n_274, n_275, n_276);
  xor g252 (n_277, n_135, n_136);
  xor g253 (n_140, n_277, n_137);
  nand g254 (n_278, n_135, n_136);
  nand g255 (n_279, n_137, n_136);
  nand g256 (n_280, n_135, n_137);
  nand g257 (n_156, n_278, n_279, n_280);
  xor g258 (n_281, n_138, n_139);
  xor g259 (n_58, n_281, n_140);
  nand g260 (n_282, n_138, n_139);
  nand g261 (n_283, n_140, n_139);
  nand g262 (n_284, n_138, n_140);
  nand g263 (n_40, n_282, n_283, n_284);
  xor g264 (n_285, in_0[5], in_1[5]);
  xor g265 (n_149, n_285, n_141);
  nand g266 (n_286, in_0[5], in_1[5]);
  nand g267 (n_287, n_141, in_1[5]);
  nand g268 (n_288, in_0[5], n_141);
  nand g269 (n_161, n_286, n_287, n_288);
  xor g270 (n_289, n_142, n_143);
  xor g271 (n_150, n_289, n_144);
  nand g272 (n_290, n_142, n_143);
  nand g273 (n_291, n_144, n_143);
  nand g274 (n_292, n_142, n_144);
  nand g275 (n_162, n_290, n_291, n_292);
  xor g276 (n_293, n_145, n_146);
  xor g277 (n_152, n_293, n_147);
  nand g278 (n_294, n_145, n_146);
  nand g279 (n_295, n_147, n_146);
  nand g280 (n_296, n_145, n_147);
  nand g281 (n_164, n_294, n_295, n_296);
  xor g282 (n_297, n_148, n_149);
  xor g283 (n_153, n_297, n_150);
  nand g284 (n_298, n_148, n_149);
  nand g285 (n_299, n_150, n_149);
  nand g286 (n_300, n_148, n_150);
  nand g287 (n_165, n_298, n_299, n_300);
  xor g288 (n_301, n_151, n_152);
  xor g289 (n_155, n_301, n_153);
  nand g290 (n_302, n_151, n_152);
  nand g291 (n_303, n_153, n_152);
  nand g292 (n_304, n_151, n_153);
  nand g293 (n_168, n_302, n_303, n_304);
  xor g294 (n_305, n_154, n_155);
  xor g295 (n_57, n_305, n_156);
  nand g296 (n_306, n_154, n_155);
  nand g297 (n_307, n_156, n_155);
  nand g298 (n_308, n_154, n_156);
  nand g299 (n_39, n_306, n_307, n_308);
  xor g300 (n_309, n_157, n_158);
  xor g301 (n_163, n_309, n_159);
  nand g302 (n_310, n_157, n_158);
  nand g303 (n_311, n_159, n_158);
  nand g304 (n_312, n_157, n_159);
  nand g305 (n_174, n_310, n_311, n_312);
  xor g306 (n_313, n_160, n_161);
  xor g307 (n_166, n_313, n_162);
  nand g308 (n_314, n_160, n_161);
  nand g309 (n_315, n_162, n_161);
  nand g310 (n_316, n_160, n_162);
  nand g311 (n_176, n_314, n_315, n_316);
  xor g312 (n_317, n_163, n_164);
  xor g313 (n_167, n_317, n_165);
  nand g314 (n_318, n_163, n_164);
  nand g315 (n_319, n_165, n_164);
  nand g316 (n_320, n_163, n_165);
  nand g317 (n_178, n_318, n_319, n_320);
  xor g318 (n_321, n_166, n_167);
  xor g319 (n_56, n_321, n_168);
  nand g320 (n_322, n_166, n_167);
  nand g321 (n_323, n_168, n_167);
  nand g322 (n_324, n_166, n_168);
  nand g323 (n_38, n_322, n_323, n_324);
  xor g324 (n_325, in_0[6], in_1[6]);
  xor g325 (n_173, n_325, n_169);
  nand g326 (n_326, in_0[6], in_1[6]);
  nand g327 (n_327, n_169, in_1[6]);
  nand g328 (n_328, in_0[6], n_169);
  nand g329 (n_182, n_326, n_327, n_328);
  xor g330 (n_329, n_170, n_171);
  xor g331 (n_175, n_329, n_172);
  nand g332 (n_330, n_170, n_171);
  nand g333 (n_331, n_172, n_171);
  nand g334 (n_332, n_170, n_172);
  nand g335 (n_181, n_330, n_331, n_332);
  xor g336 (n_333, n_173, n_174);
  xor g337 (n_177, n_333, n_175);
  nand g338 (n_334, n_173, n_174);
  nand g339 (n_335, n_175, n_174);
  nand g340 (n_336, n_173, n_175);
  nand g341 (n_184, n_334, n_335, n_336);
  xor g342 (n_337, n_176, n_177);
  xor g343 (n_55, n_337, n_178);
  nand g344 (n_338, n_176, n_177);
  nand g345 (n_339, n_178, n_177);
  nand g346 (n_340, n_176, n_178);
  nand g347 (n_54, n_338, n_339, n_340);
  xor g348 (n_341, n_179, n_180);
  xor g349 (n_183, n_341, n_181);
  nand g350 (n_342, n_179, n_180);
  nand g351 (n_343, n_181, n_180);
  nand g352 (n_344, n_179, n_181);
  nand g353 (n_188, n_342, n_343, n_344);
  xor g354 (n_345, n_182, n_183);
  xor g355 (n_37, n_345, n_184);
  nand g356 (n_346, n_182, n_183);
  nand g357 (n_347, n_184, n_183);
  nand g358 (n_348, n_182, n_184);
  nand g359 (n_53, n_346, n_347, n_348);
  xor g360 (n_349, in_0[7], in_1[7]);
  xor g361 (n_187, n_349, n_185);
  nand g362 (n_350, in_0[7], in_1[7]);
  nand g363 (n_351, n_185, in_1[7]);
  nand g364 (n_352, in_0[7], n_185);
  nand g365 (n_35, n_350, n_351, n_352);
  xor g366 (n_353, n_186, n_187);
  xor g367 (n_36, n_353, n_188);
  nand g368 (n_354, n_186, n_187);
  nand g369 (n_355, n_188, n_187);
  nand g370 (n_356, n_186, n_188);
  nand g371 (n_52, n_354, n_355, n_356);
  nand g374 (n_358, in_1[0], in_0[0]);
  nor g379 (n_370, n_48, n_65);
  nand g380 (n_365, n_48, n_65);
  nor g381 (n_366, n_47, n_64);
  nand g382 (n_367, n_47, n_64);
  nor g383 (n_376, n_46, n_63);
  nand g384 (n_371, n_46, n_63);
  nor g385 (n_372, n_45, n_62);
  nand g386 (n_373, n_45, n_62);
  nor g387 (n_382, n_44, n_61);
  nand g388 (n_377, n_44, n_61);
  nor g389 (n_378, n_43, n_60);
  nand g390 (n_379, n_43, n_60);
  nor g391 (n_388, n_42, n_59);
  nand g392 (n_383, n_42, n_59);
  nor g393 (n_384, n_41, n_58);
  nand g394 (n_385, n_41, n_58);
  nor g395 (n_394, n_40, n_57);
  nand g396 (n_389, n_40, n_57);
  nor g397 (n_390, n_39, n_56);
  nand g398 (n_391, n_39, n_56);
  nor g399 (n_400, n_38, n_55);
  nand g400 (n_395, n_38, n_55);
  nor g401 (n_396, n_37, n_54);
  nand g402 (n_397, n_37, n_54);
  nor g403 (n_406, n_36, n_53);
  nand g404 (n_401, n_36, n_53);
  nor g405 (n_402, n_35, n_52);
  nand g406 (n_403, n_35, n_52);
  nor g412 (n_368, n_365, n_366);
  nor g416 (n_374, n_371, n_372);
  nor g419 (n_416, n_376, n_372);
  nor g420 (n_380, n_377, n_378);
  nor g423 (n_418, n_382, n_378);
  nor g424 (n_386, n_383, n_384);
  nor g427 (n_426, n_388, n_384);
  nor g57 (n_392, n_389, n_390);
  nor g60 (n_428, n_394, n_390);
  nor g61 (n_398, n_395, n_396);
  nor g64 (n_436, n_400, n_396);
  nor g65 (n_404, n_401, n_402);
  nor g68 (n_438, n_406, n_402);
  nor g74 (n_414, n_382, n_413);
  nand g83 (n_451, n_416, n_418);
  nor g84 (n_424, n_394, n_423);
  nand g93 (n_458, n_426, n_428);
  nor g94 (n_434, n_406, n_433);
  nand g103 (n_466, n_436, n_438);
  nand g428 (n_503, n_371, n_543);
  nand g430 (n_505, n_413, n_544);
  nand g433 (n_508, n_550, n_551);
  nand g436 (n_470, n_561, n_562);
  nor g437 (n_456, n_400, n_455);
  nor g440 (n_480, n_400, n_458);
  nor g446 (n_464, n_462, n_455);
  nor g449 (n_486, n_458, n_462);
  nor g450 (n_468, n_466, n_455);
  nor g453 (n_489, n_458, n_466);
  nand g456 (n_512, n_383, n_572);
  nand g457 (n_473, n_426, n_470);
  nand g458 (n_514, n_423, n_473);
  nand g461 (n_517, n_566, n_573);
  nand g464 (n_520, n_455, n_574);
  nand g465 (n_482, n_480, n_470);
  nand g466 (n_523, n_576, n_482);
  nand g467 (n_485, n_569, n_470);
  nand g468 (n_525, n_577, n_485);
  nand g469 (n_488, n_486, n_470);
  nand g470 (n_528, n_578, n_488);
  nand g471 (n_491, n_489, n_470);
  nand g472 (out_0[16], n_579, n_491);
  xnor g485 (out_0[5], n_503, n_546);
  xnor g487 (out_0[6], n_505, n_547);
  xnor g490 (out_0[7], n_508, n_552);
  xnor g492 (out_0[8], n_470, n_553);
  xnor g495 (out_0[9], n_512, n_558);
  xnor g497 (out_0[10], n_514, n_559);
  xnor g500 (out_0[11], n_517, n_563);
  xnor g503 (out_0[12], n_520, n_564);
  xnor g506 (out_0[13], n_523, n_565);
  xnor g508 (out_0[14], n_525, n_554);
  xnor g511 (out_0[15], n_528, n_555);
  xor g514 (out_0[0], in_0[0], in_1[0]);
  not g515 (out_0[1], n_358);
  or g516 (n_535, wc, n_370);
  not gc (wc, n_365);
  and g517 (n_536, wc0, n_367);
  not gc0 (wc0, n_368);
  not g519 (out_0[2], n_535);
  or g520 (n_539, wc1, n_366);
  not gc1 (wc1, n_367);
  or g521 (n_540, wc2, n_376);
  not gc2 (wc2, n_371);
  xor g523 (out_0[3], n_365, n_539);
  and g524 (n_413, wc3, n_373);
  not gc3 (wc3, n_374);
  or g525 (n_542, wc4, n_382);
  not gc4 (wc4, n_416);
  or g526 (n_543, n_376, n_536);
  or g527 (n_544, n_536, wc5);
  not gc5 (wc5, n_416);
  xor g528 (out_0[4], n_536, n_540);
  or g529 (n_546, wc6, n_372);
  not gc6 (wc6, n_373);
  or g530 (n_547, wc7, n_382);
  not gc7 (wc7, n_377);
  and g531 (n_548, wc8, n_379);
  not gc8 (wc8, n_380);
  and g532 (n_549, wc9, n_403);
  not gc9 (wc9, n_404);
  and g533 (n_550, wc10, n_377);
  not gc10 (wc10, n_414);
  or g534 (n_551, n_536, n_542);
  or g535 (n_552, wc11, n_378);
  not gc11 (wc11, n_379);
  or g536 (n_553, wc12, n_388);
  not gc12 (wc12, n_383);
  or g537 (n_554, wc13, n_406);
  not gc13 (wc13, n_401);
  or g538 (n_555, wc14, n_402);
  not gc14 (wc14, n_403);
  and g539 (n_423, wc15, n_385);
  not gc15 (wc15, n_386);
  and g540 (n_556, wc16, n_418);
  not gc16 (wc16, n_413);
  or g541 (n_557, wc17, n_394);
  not gc17 (wc17, n_426);
  or g542 (n_558, wc18, n_384);
  not gc18 (wc18, n_385);
  or g543 (n_559, wc19, n_394);
  not gc19 (wc19, n_389);
  and g544 (n_560, wc20, n_391);
  not gc20 (wc20, n_392);
  and g545 (n_433, wc21, n_397);
  not gc21 (wc21, n_398);
  and g546 (n_561, wc22, n_548);
  not gc22 (wc22, n_556);
  or g547 (n_462, wc23, n_406);
  not gc23 (wc23, n_436);
  or g548 (n_562, n_451, n_536);
  or g549 (n_563, wc24, n_390);
  not gc24 (wc24, n_391);
  or g550 (n_564, wc25, n_400);
  not gc25 (wc25, n_395);
  or g551 (n_565, wc26, n_396);
  not gc26 (wc26, n_397);
  and g552 (n_566, wc27, n_389);
  not gc27 (wc27, n_424);
  and g553 (n_567, wc28, n_428);
  not gc28 (wc28, n_423);
  and g554 (n_568, wc29, n_438);
  not gc29 (wc29, n_433);
  and g555 (n_569, wc30, n_436);
  not gc30 (wc30, n_458);
  and g556 (n_455, wc31, n_560);
  not gc31 (wc31, n_567);
  and g557 (n_570, wc32, n_401);
  not gc32 (wc32, n_434);
  and g558 (n_571, wc33, n_549);
  not gc33 (wc33, n_568);
  or g559 (n_572, wc34, n_388);
  not gc34 (wc34, n_470);
  or g560 (n_573, n_557, wc35);
  not gc35 (wc35, n_470);
  or g561 (n_574, wc36, n_458);
  not gc36 (wc36, n_470);
  and g562 (n_575, wc37, n_436);
  not gc37 (wc37, n_455);
  and g563 (n_576, wc38, n_395);
  not gc38 (wc38, n_456);
  and g564 (n_577, wc39, n_433);
  not gc39 (wc39, n_575);
  and g565 (n_578, n_570, wc40);
  not gc40 (wc40, n_464);
  and g566 (n_579, n_571, wc41);
  not gc41 (wc41, n_468);
endmodule

module csa_tree_distance1_add1033_group_329_GENERIC(in_0, in_1, out_0);
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  csa_tree_distance1_add1033_group_329_GENERIC_REAL g1(.in_0 (in_0),
       .in_1 (in_1), .out_0 (out_0));
endmodule

module csa_tree_distance2_add1032_group_331_GENERIC_REAL(in_0, in_1,
     out_0);
// synthesis_equation "assign out_0 = ( ( in_0 * in_0 )  + ( in_1 * in_1 )  )  ;"
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_358, n_365, n_366, n_367, n_368, n_370;
  wire n_371, n_372, n_373, n_374, n_376, n_377, n_378, n_379;
  wire n_380, n_382, n_383, n_384, n_385, n_386, n_388, n_389;
  wire n_390, n_391, n_392, n_394, n_395, n_396, n_397, n_398;
  wire n_400, n_401, n_402, n_403, n_404, n_406, n_413, n_414;
  wire n_416, n_418, n_423, n_424, n_426, n_428, n_433, n_434;
  wire n_436, n_438, n_451, n_455, n_456, n_458, n_462, n_464;
  wire n_466, n_468, n_470, n_473, n_480, n_482, n_485, n_486;
  wire n_488, n_489, n_491, n_503, n_505, n_508, n_512, n_514;
  wire n_517, n_520, n_523, n_525, n_528, n_535, n_536, n_539;
  wire n_540, n_542, n_543, n_544, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579;
  and g1 (n_48, in_0[0], in_0[1]);
  and g2 (n_70, in_0[0], in_0[2]);
  and g3 (n_74, in_0[1], in_0[2]);
  and g4 (n_75, in_0[0], in_0[3]);
  and g5 (n_78, in_0[1], in_0[3]);
  and g6 (n_86, in_0[2], in_0[3]);
  and g7 (n_79, in_0[0], in_0[4]);
  and g8 (n_90, in_0[1], in_0[4]);
  and g9 (n_98, in_0[2], in_0[4]);
  and g10 (n_109, in_0[3], in_0[4]);
  and g11 (n_87, in_0[0], in_0[5]);
  and g12 (n_99, in_0[1], in_0[5]);
  and g13 (n_67, in_0[2], in_0[5]);
  and g14 (n_124, in_0[3], in_0[5]);
  and g15 (n_141, in_0[4], in_0[5]);
  and g16 (n_50, in_0[0], in_0[6]);
  and g17 (n_110, in_0[1], in_0[6]);
  and g18 (n_125, in_0[2], in_0[6]);
  and g19 (n_145, in_0[3], in_0[6]);
  and g20 (n_157, in_0[4], in_0[6]);
  and g21 (n_170, in_0[5], in_0[6]);
  and g22 (n_113, in_0[0], in_0[7]);
  and g23 (n_128, in_0[1], in_0[7]);
  and g24 (n_142, in_0[2], in_0[7]);
  and g25 (n_158, in_0[3], in_0[7]);
  and g26 (n_171, in_0[4], in_0[7]);
  and g27 (n_179, in_0[5], in_0[7]);
  and g28 (n_185, in_0[6], in_0[7]);
  and g29 (n_69, in_1[0], in_1[1]);
  and g30 (n_71, in_1[0], in_1[2]);
  and g31 (n_73, in_1[1], in_1[2]);
  and g32 (n_72, in_1[0], in_1[3]);
  and g33 (n_81, in_1[1], in_1[3]);
  and g34 (n_89, in_1[2], in_1[3]);
  and g35 (n_80, in_1[0], in_1[4]);
  and g36 (n_91, in_1[1], in_1[4]);
  and g37 (n_100, in_1[2], in_1[4]);
  and g38 (n_66, in_1[3], in_1[4]);
  and g39 (n_88, in_1[0], in_1[5]);
  and g40 (n_49, in_1[1], in_1[5]);
  and g41 (n_111, in_1[2], in_1[5]);
  and g42 (n_126, in_1[3], in_1[5]);
  and g43 (n_144, in_1[4], in_1[5]);
  and g44 (n_51, in_1[0], in_1[6]);
  and g45 (n_112, in_1[1], in_1[6]);
  and g46 (n_127, in_1[2], in_1[6]);
  and g47 (n_146, in_1[3], in_1[6]);
  and g48 (n_160, in_1[4], in_1[6]);
  and g49 (n_169, in_1[5], in_1[6]);
  and g50 (n_114, in_1[0], in_1[7]);
  and g51 (n_129, in_1[1], in_1[7]);
  and g52 (n_143, in_1[2], in_1[7]);
  and g53 (n_159, in_1[3], in_1[7]);
  and g54 (n_172, in_1[4], in_1[7]);
  and g55 (n_180, in_1[5], in_1[7]);
  and g56 (n_186, in_1[6], in_1[7]);
  xor g106 (n_189, in_0[1], in_1[1]);
  xor g107 (n_65, n_189, n_69);
  nand g108 (n_190, in_0[1], in_1[1]);
  nand g109 (n_191, n_69, in_1[1]);
  nand g110 (n_192, in_0[1], n_69);
  nand g111 (n_64, n_190, n_191, n_192);
  xor g112 (n_47, n_70, n_71);
  and g113 (n_77, n_70, n_71);
  xor g114 (n_76, in_0[2], in_1[2]);
  and g115 (n_82, in_0[2], in_1[2]);
  xor g116 (n_193, n_72, n_73);
  xor g117 (n_46, n_193, n_74);
  nand g118 (n_194, n_72, n_73);
  nand g119 (n_195, n_74, n_73);
  nand g120 (n_196, n_72, n_74);
  nand g121 (n_84, n_194, n_195, n_196);
  xor g122 (n_197, n_75, n_76);
  xor g123 (n_63, n_197, n_77);
  nand g124 (n_198, n_75, n_76);
  nand g125 (n_199, n_77, n_76);
  nand g126 (n_200, n_75, n_77);
  nand g127 (n_45, n_198, n_199, n_200);
  xor g128 (n_83, n_78, n_79);
  and g129 (n_93, n_78, n_79);
  xor g130 (n_201, n_80, n_81);
  xor g131 (n_85, n_201, n_82);
  nand g132 (n_202, n_80, n_81);
  nand g133 (n_203, n_82, n_81);
  nand g134 (n_204, n_80, n_82);
  nand g135 (n_95, n_202, n_203, n_204);
  xor g136 (n_205, n_83, n_84);
  xor g137 (n_62, n_205, n_85);
  nand g138 (n_206, n_83, n_84);
  nand g139 (n_207, n_85, n_84);
  nand g140 (n_208, n_83, n_85);
  nand g141 (n_44, n_206, n_207, n_208);
  xor g142 (n_92, in_0[3], in_1[3]);
  and g143 (n_101, in_0[3], in_1[3]);
  xor g144 (n_209, n_86, n_87);
  xor g145 (n_96, n_209, n_88);
  nand g146 (n_210, n_86, n_87);
  nand g147 (n_211, n_88, n_87);
  nand g148 (n_212, n_86, n_88);
  nand g149 (n_103, n_210, n_211, n_212);
  xor g150 (n_213, n_89, n_90);
  xor g151 (n_94, n_213, n_91);
  nand g152 (n_214, n_89, n_90);
  nand g153 (n_215, n_91, n_90);
  nand g154 (n_216, n_89, n_91);
  nand g155 (n_104, n_214, n_215, n_216);
  xor g156 (n_217, n_92, n_93);
  xor g157 (n_97, n_217, n_94);
  nand g158 (n_218, n_92, n_93);
  nand g159 (n_219, n_94, n_93);
  nand g160 (n_220, n_92, n_94);
  nand g161 (n_108, n_218, n_219, n_220);
  xor g162 (n_221, n_95, n_96);
  xor g163 (n_61, n_221, n_97);
  nand g164 (n_222, n_95, n_96);
  nand g165 (n_223, n_97, n_96);
  nand g166 (n_224, n_95, n_97);
  nand g167 (n_43, n_222, n_223, n_224);
  xor g168 (n_102, n_98, n_99);
  and g169 (n_115, n_98, n_99);
  xor g170 (n_225, n_100, n_49);
  xor g171 (n_105, n_225, n_50);
  nand g172 (n_226, n_100, n_49);
  nand g173 (n_227, n_50, n_49);
  nand g174 (n_228, n_100, n_50);
  nand g175 (n_116, n_226, n_227, n_228);
  xor g176 (n_229, n_51, n_101);
  xor g177 (n_106, n_229, n_102);
  nand g178 (n_230, n_51, n_101);
  nand g179 (n_231, n_102, n_101);
  nand g180 (n_232, n_51, n_102);
  nand g181 (n_120, n_230, n_231, n_232);
  xor g182 (n_233, n_103, n_104);
  xor g183 (n_107, n_233, n_105);
  nand g184 (n_234, n_103, n_104);
  nand g185 (n_235, n_105, n_104);
  nand g186 (n_236, n_103, n_105);
  nand g187 (n_121, n_234, n_235, n_236);
  xor g188 (n_237, n_106, n_107);
  xor g189 (n_60, n_237, n_108);
  nand g190 (n_238, n_106, n_107);
  nand g191 (n_239, n_108, n_107);
  nand g192 (n_240, n_106, n_108);
  nand g193 (n_42, n_238, n_239, n_240);
  xor g194 (n_68, in_0[4], in_1[4]);
  and g195 (n_130, in_0[4], in_1[4]);
  xor g196 (n_241, n_109, n_110);
  xor g197 (n_117, n_241, n_111);
  nand g198 (n_242, n_109, n_110);
  nand g199 (n_243, n_111, n_110);
  nand g200 (n_244, n_109, n_111);
  nand g201 (n_133, n_242, n_243, n_244);
  xor g202 (n_245, n_112, n_113);
  xor g203 (n_119, n_245, n_114);
  nand g204 (n_246, n_112, n_113);
  nand g205 (n_247, n_114, n_113);
  nand g206 (n_248, n_112, n_114);
  nand g207 (n_132, n_246, n_247, n_248);
  xor g208 (n_249, n_66, n_67);
  xor g209 (n_118, n_249, n_68);
  nand g210 (n_250, n_66, n_67);
  nand g211 (n_251, n_68, n_67);
  nand g212 (n_252, n_66, n_68);
  nand g213 (n_134, n_250, n_251, n_252);
  xor g214 (n_253, n_115, n_116);
  xor g215 (n_122, n_253, n_117);
  nand g216 (n_254, n_115, n_116);
  nand g217 (n_255, n_117, n_116);
  nand g218 (n_256, n_115, n_117);
  nand g219 (n_138, n_254, n_255, n_256);
  xor g220 (n_257, n_118, n_119);
  xor g221 (n_123, n_257, n_120);
  nand g222 (n_258, n_118, n_119);
  nand g223 (n_259, n_120, n_119);
  nand g224 (n_260, n_118, n_120);
  nand g225 (n_139, n_258, n_259, n_260);
  xor g226 (n_261, n_121, n_122);
  xor g227 (n_59, n_261, n_123);
  nand g228 (n_262, n_121, n_122);
  nand g229 (n_263, n_123, n_122);
  nand g230 (n_264, n_121, n_123);
  nand g231 (n_41, n_262, n_263, n_264);
  xor g232 (n_131, n_124, n_125);
  and g233 (n_147, n_124, n_125);
  xor g234 (n_265, n_126, n_127);
  xor g235 (n_135, n_265, n_128);
  nand g236 (n_266, n_126, n_127);
  nand g237 (n_267, n_128, n_127);
  nand g238 (n_268, n_126, n_128);
  nand g239 (n_148, n_266, n_267, n_268);
  xor g240 (n_269, n_129, n_130);
  xor g241 (n_136, n_269, n_131);
  nand g242 (n_270, n_129, n_130);
  nand g243 (n_271, n_131, n_130);
  nand g244 (n_272, n_129, n_131);
  nand g245 (n_151, n_270, n_271, n_272);
  xor g246 (n_273, n_132, n_133);
  xor g247 (n_137, n_273, n_134);
  nand g248 (n_274, n_132, n_133);
  nand g249 (n_275, n_134, n_133);
  nand g250 (n_276, n_132, n_134);
  nand g251 (n_154, n_274, n_275, n_276);
  xor g252 (n_277, n_135, n_136);
  xor g253 (n_140, n_277, n_137);
  nand g254 (n_278, n_135, n_136);
  nand g255 (n_279, n_137, n_136);
  nand g256 (n_280, n_135, n_137);
  nand g257 (n_156, n_278, n_279, n_280);
  xor g258 (n_281, n_138, n_139);
  xor g259 (n_58, n_281, n_140);
  nand g260 (n_282, n_138, n_139);
  nand g261 (n_283, n_140, n_139);
  nand g262 (n_284, n_138, n_140);
  nand g263 (n_40, n_282, n_283, n_284);
  xor g264 (n_285, in_0[5], in_1[5]);
  xor g265 (n_149, n_285, n_141);
  nand g266 (n_286, in_0[5], in_1[5]);
  nand g267 (n_287, n_141, in_1[5]);
  nand g268 (n_288, in_0[5], n_141);
  nand g269 (n_161, n_286, n_287, n_288);
  xor g270 (n_289, n_142, n_143);
  xor g271 (n_150, n_289, n_144);
  nand g272 (n_290, n_142, n_143);
  nand g273 (n_291, n_144, n_143);
  nand g274 (n_292, n_142, n_144);
  nand g275 (n_162, n_290, n_291, n_292);
  xor g276 (n_293, n_145, n_146);
  xor g277 (n_152, n_293, n_147);
  nand g278 (n_294, n_145, n_146);
  nand g279 (n_295, n_147, n_146);
  nand g280 (n_296, n_145, n_147);
  nand g281 (n_164, n_294, n_295, n_296);
  xor g282 (n_297, n_148, n_149);
  xor g283 (n_153, n_297, n_150);
  nand g284 (n_298, n_148, n_149);
  nand g285 (n_299, n_150, n_149);
  nand g286 (n_300, n_148, n_150);
  nand g287 (n_165, n_298, n_299, n_300);
  xor g288 (n_301, n_151, n_152);
  xor g289 (n_155, n_301, n_153);
  nand g290 (n_302, n_151, n_152);
  nand g291 (n_303, n_153, n_152);
  nand g292 (n_304, n_151, n_153);
  nand g293 (n_168, n_302, n_303, n_304);
  xor g294 (n_305, n_154, n_155);
  xor g295 (n_57, n_305, n_156);
  nand g296 (n_306, n_154, n_155);
  nand g297 (n_307, n_156, n_155);
  nand g298 (n_308, n_154, n_156);
  nand g299 (n_39, n_306, n_307, n_308);
  xor g300 (n_309, n_157, n_158);
  xor g301 (n_163, n_309, n_159);
  nand g302 (n_310, n_157, n_158);
  nand g303 (n_311, n_159, n_158);
  nand g304 (n_312, n_157, n_159);
  nand g305 (n_174, n_310, n_311, n_312);
  xor g306 (n_313, n_160, n_161);
  xor g307 (n_166, n_313, n_162);
  nand g308 (n_314, n_160, n_161);
  nand g309 (n_315, n_162, n_161);
  nand g310 (n_316, n_160, n_162);
  nand g311 (n_176, n_314, n_315, n_316);
  xor g312 (n_317, n_163, n_164);
  xor g313 (n_167, n_317, n_165);
  nand g314 (n_318, n_163, n_164);
  nand g315 (n_319, n_165, n_164);
  nand g316 (n_320, n_163, n_165);
  nand g317 (n_178, n_318, n_319, n_320);
  xor g318 (n_321, n_166, n_167);
  xor g319 (n_56, n_321, n_168);
  nand g320 (n_322, n_166, n_167);
  nand g321 (n_323, n_168, n_167);
  nand g322 (n_324, n_166, n_168);
  nand g323 (n_38, n_322, n_323, n_324);
  xor g324 (n_325, in_0[6], in_1[6]);
  xor g325 (n_173, n_325, n_169);
  nand g326 (n_326, in_0[6], in_1[6]);
  nand g327 (n_327, n_169, in_1[6]);
  nand g328 (n_328, in_0[6], n_169);
  nand g329 (n_182, n_326, n_327, n_328);
  xor g330 (n_329, n_170, n_171);
  xor g331 (n_175, n_329, n_172);
  nand g332 (n_330, n_170, n_171);
  nand g333 (n_331, n_172, n_171);
  nand g334 (n_332, n_170, n_172);
  nand g335 (n_181, n_330, n_331, n_332);
  xor g336 (n_333, n_173, n_174);
  xor g337 (n_177, n_333, n_175);
  nand g338 (n_334, n_173, n_174);
  nand g339 (n_335, n_175, n_174);
  nand g340 (n_336, n_173, n_175);
  nand g341 (n_184, n_334, n_335, n_336);
  xor g342 (n_337, n_176, n_177);
  xor g343 (n_55, n_337, n_178);
  nand g344 (n_338, n_176, n_177);
  nand g345 (n_339, n_178, n_177);
  nand g346 (n_340, n_176, n_178);
  nand g347 (n_54, n_338, n_339, n_340);
  xor g348 (n_341, n_179, n_180);
  xor g349 (n_183, n_341, n_181);
  nand g350 (n_342, n_179, n_180);
  nand g351 (n_343, n_181, n_180);
  nand g352 (n_344, n_179, n_181);
  nand g353 (n_188, n_342, n_343, n_344);
  xor g354 (n_345, n_182, n_183);
  xor g355 (n_37, n_345, n_184);
  nand g356 (n_346, n_182, n_183);
  nand g357 (n_347, n_184, n_183);
  nand g358 (n_348, n_182, n_184);
  nand g359 (n_53, n_346, n_347, n_348);
  xor g360 (n_349, in_0[7], in_1[7]);
  xor g361 (n_187, n_349, n_185);
  nand g362 (n_350, in_0[7], in_1[7]);
  nand g363 (n_351, n_185, in_1[7]);
  nand g364 (n_352, in_0[7], n_185);
  nand g365 (n_35, n_350, n_351, n_352);
  xor g366 (n_353, n_186, n_187);
  xor g367 (n_36, n_353, n_188);
  nand g368 (n_354, n_186, n_187);
  nand g369 (n_355, n_188, n_187);
  nand g370 (n_356, n_186, n_188);
  nand g371 (n_52, n_354, n_355, n_356);
  nand g374 (n_358, in_1[0], in_0[0]);
  nor g379 (n_370, n_48, n_65);
  nand g380 (n_365, n_48, n_65);
  nor g381 (n_366, n_47, n_64);
  nand g382 (n_367, n_47, n_64);
  nor g383 (n_376, n_46, n_63);
  nand g384 (n_371, n_46, n_63);
  nor g385 (n_372, n_45, n_62);
  nand g386 (n_373, n_45, n_62);
  nor g387 (n_382, n_44, n_61);
  nand g388 (n_377, n_44, n_61);
  nor g389 (n_378, n_43, n_60);
  nand g390 (n_379, n_43, n_60);
  nor g391 (n_388, n_42, n_59);
  nand g392 (n_383, n_42, n_59);
  nor g393 (n_384, n_41, n_58);
  nand g394 (n_385, n_41, n_58);
  nor g395 (n_394, n_40, n_57);
  nand g396 (n_389, n_40, n_57);
  nor g397 (n_390, n_39, n_56);
  nand g398 (n_391, n_39, n_56);
  nor g399 (n_400, n_38, n_55);
  nand g400 (n_395, n_38, n_55);
  nor g401 (n_396, n_37, n_54);
  nand g402 (n_397, n_37, n_54);
  nor g403 (n_406, n_36, n_53);
  nand g404 (n_401, n_36, n_53);
  nor g405 (n_402, n_35, n_52);
  nand g406 (n_403, n_35, n_52);
  nor g412 (n_368, n_365, n_366);
  nor g416 (n_374, n_371, n_372);
  nor g419 (n_416, n_376, n_372);
  nor g420 (n_380, n_377, n_378);
  nor g423 (n_418, n_382, n_378);
  nor g424 (n_386, n_383, n_384);
  nor g427 (n_426, n_388, n_384);
  nor g57 (n_392, n_389, n_390);
  nor g60 (n_428, n_394, n_390);
  nor g61 (n_398, n_395, n_396);
  nor g64 (n_436, n_400, n_396);
  nor g65 (n_404, n_401, n_402);
  nor g68 (n_438, n_406, n_402);
  nor g74 (n_414, n_382, n_413);
  nand g83 (n_451, n_416, n_418);
  nor g84 (n_424, n_394, n_423);
  nand g93 (n_458, n_426, n_428);
  nor g94 (n_434, n_406, n_433);
  nand g103 (n_466, n_436, n_438);
  nand g428 (n_503, n_371, n_543);
  nand g430 (n_505, n_413, n_544);
  nand g433 (n_508, n_550, n_551);
  nand g436 (n_470, n_561, n_562);
  nor g437 (n_456, n_400, n_455);
  nor g440 (n_480, n_400, n_458);
  nor g446 (n_464, n_462, n_455);
  nor g449 (n_486, n_458, n_462);
  nor g450 (n_468, n_466, n_455);
  nor g453 (n_489, n_458, n_466);
  nand g456 (n_512, n_383, n_572);
  nand g457 (n_473, n_426, n_470);
  nand g458 (n_514, n_423, n_473);
  nand g461 (n_517, n_566, n_573);
  nand g464 (n_520, n_455, n_574);
  nand g465 (n_482, n_480, n_470);
  nand g466 (n_523, n_576, n_482);
  nand g467 (n_485, n_569, n_470);
  nand g468 (n_525, n_577, n_485);
  nand g469 (n_488, n_486, n_470);
  nand g470 (n_528, n_578, n_488);
  nand g471 (n_491, n_489, n_470);
  nand g472 (out_0[16], n_579, n_491);
  xnor g485 (out_0[5], n_503, n_546);
  xnor g487 (out_0[6], n_505, n_547);
  xnor g490 (out_0[7], n_508, n_552);
  xnor g492 (out_0[8], n_470, n_553);
  xnor g495 (out_0[9], n_512, n_558);
  xnor g497 (out_0[10], n_514, n_559);
  xnor g500 (out_0[11], n_517, n_563);
  xnor g503 (out_0[12], n_520, n_564);
  xnor g506 (out_0[13], n_523, n_565);
  xnor g508 (out_0[14], n_525, n_554);
  xnor g511 (out_0[15], n_528, n_555);
  xor g514 (out_0[0], in_0[0], in_1[0]);
  not g515 (out_0[1], n_358);
  or g516 (n_535, wc, n_370);
  not gc (wc, n_365);
  and g517 (n_536, wc0, n_367);
  not gc0 (wc0, n_368);
  not g519 (out_0[2], n_535);
  or g520 (n_539, wc1, n_366);
  not gc1 (wc1, n_367);
  or g521 (n_540, wc2, n_376);
  not gc2 (wc2, n_371);
  xor g523 (out_0[3], n_365, n_539);
  and g524 (n_413, wc3, n_373);
  not gc3 (wc3, n_374);
  or g525 (n_542, wc4, n_382);
  not gc4 (wc4, n_416);
  or g526 (n_543, n_376, n_536);
  or g527 (n_544, n_536, wc5);
  not gc5 (wc5, n_416);
  xor g528 (out_0[4], n_536, n_540);
  or g529 (n_546, wc6, n_372);
  not gc6 (wc6, n_373);
  or g530 (n_547, wc7, n_382);
  not gc7 (wc7, n_377);
  and g531 (n_548, wc8, n_379);
  not gc8 (wc8, n_380);
  and g532 (n_549, wc9, n_403);
  not gc9 (wc9, n_404);
  and g533 (n_550, wc10, n_377);
  not gc10 (wc10, n_414);
  or g534 (n_551, n_536, n_542);
  or g535 (n_552, wc11, n_378);
  not gc11 (wc11, n_379);
  or g536 (n_553, wc12, n_388);
  not gc12 (wc12, n_383);
  or g537 (n_554, wc13, n_406);
  not gc13 (wc13, n_401);
  or g538 (n_555, wc14, n_402);
  not gc14 (wc14, n_403);
  and g539 (n_423, wc15, n_385);
  not gc15 (wc15, n_386);
  and g540 (n_556, wc16, n_418);
  not gc16 (wc16, n_413);
  or g541 (n_557, wc17, n_394);
  not gc17 (wc17, n_426);
  or g542 (n_558, wc18, n_384);
  not gc18 (wc18, n_385);
  or g543 (n_559, wc19, n_394);
  not gc19 (wc19, n_389);
  and g544 (n_560, wc20, n_391);
  not gc20 (wc20, n_392);
  and g545 (n_433, wc21, n_397);
  not gc21 (wc21, n_398);
  and g546 (n_561, wc22, n_548);
  not gc22 (wc22, n_556);
  or g547 (n_462, wc23, n_406);
  not gc23 (wc23, n_436);
  or g548 (n_562, n_451, n_536);
  or g549 (n_563, wc24, n_390);
  not gc24 (wc24, n_391);
  or g550 (n_564, wc25, n_400);
  not gc25 (wc25, n_395);
  or g551 (n_565, wc26, n_396);
  not gc26 (wc26, n_397);
  and g552 (n_566, wc27, n_389);
  not gc27 (wc27, n_424);
  and g553 (n_567, wc28, n_428);
  not gc28 (wc28, n_423);
  and g554 (n_568, wc29, n_438);
  not gc29 (wc29, n_433);
  and g555 (n_569, wc30, n_436);
  not gc30 (wc30, n_458);
  and g556 (n_455, wc31, n_560);
  not gc31 (wc31, n_567);
  and g557 (n_570, wc32, n_401);
  not gc32 (wc32, n_434);
  and g558 (n_571, wc33, n_549);
  not gc33 (wc33, n_568);
  or g559 (n_572, wc34, n_388);
  not gc34 (wc34, n_470);
  or g560 (n_573, n_557, wc35);
  not gc35 (wc35, n_470);
  or g561 (n_574, wc36, n_458);
  not gc36 (wc36, n_470);
  and g562 (n_575, wc37, n_436);
  not gc37 (wc37, n_455);
  and g563 (n_576, wc38, n_395);
  not gc38 (wc38, n_456);
  and g564 (n_577, wc39, n_433);
  not gc39 (wc39, n_575);
  and g565 (n_578, n_570, wc40);
  not gc40 (wc40, n_464);
  and g566 (n_579, n_571, wc41);
  not gc41 (wc41, n_468);
endmodule

module csa_tree_distance2_add1032_group_331_GENERIC(in_0, in_1, out_0);
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  csa_tree_distance2_add1032_group_331_GENERIC_REAL g1(.in_0 (in_0),
       .in_1 (in_1), .out_0 (out_0));
endmodule

module csa_tree_distance3_add1031_group_333_GENERIC_REAL(in_0, in_1,
     out_0);
// synthesis_equation "assign out_0 = ( ( in_0 * in_0 )  + ( in_1 * in_1 )  )  ;"
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_358, n_365, n_366, n_367, n_368, n_370;
  wire n_371, n_372, n_373, n_374, n_376, n_377, n_378, n_379;
  wire n_380, n_382, n_383, n_384, n_385, n_386, n_388, n_389;
  wire n_390, n_391, n_392, n_394, n_395, n_396, n_397, n_398;
  wire n_400, n_401, n_402, n_403, n_404, n_406, n_413, n_414;
  wire n_416, n_418, n_423, n_424, n_426, n_428, n_433, n_434;
  wire n_436, n_438, n_451, n_455, n_456, n_458, n_462, n_464;
  wire n_466, n_468, n_470, n_473, n_480, n_482, n_485, n_486;
  wire n_488, n_489, n_491, n_503, n_505, n_508, n_512, n_514;
  wire n_517, n_520, n_523, n_525, n_528, n_535, n_536, n_539;
  wire n_540, n_542, n_543, n_544, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579;
  and g1 (n_48, in_0[0], in_0[1]);
  and g2 (n_70, in_0[0], in_0[2]);
  and g3 (n_74, in_0[1], in_0[2]);
  and g4 (n_75, in_0[0], in_0[3]);
  and g5 (n_78, in_0[1], in_0[3]);
  and g6 (n_86, in_0[2], in_0[3]);
  and g7 (n_79, in_0[0], in_0[4]);
  and g8 (n_90, in_0[1], in_0[4]);
  and g9 (n_98, in_0[2], in_0[4]);
  and g10 (n_109, in_0[3], in_0[4]);
  and g11 (n_87, in_0[0], in_0[5]);
  and g12 (n_99, in_0[1], in_0[5]);
  and g13 (n_67, in_0[2], in_0[5]);
  and g14 (n_124, in_0[3], in_0[5]);
  and g15 (n_141, in_0[4], in_0[5]);
  and g16 (n_50, in_0[0], in_0[6]);
  and g17 (n_110, in_0[1], in_0[6]);
  and g18 (n_125, in_0[2], in_0[6]);
  and g19 (n_145, in_0[3], in_0[6]);
  and g20 (n_157, in_0[4], in_0[6]);
  and g21 (n_170, in_0[5], in_0[6]);
  and g22 (n_113, in_0[0], in_0[7]);
  and g23 (n_128, in_0[1], in_0[7]);
  and g24 (n_142, in_0[2], in_0[7]);
  and g25 (n_158, in_0[3], in_0[7]);
  and g26 (n_171, in_0[4], in_0[7]);
  and g27 (n_179, in_0[5], in_0[7]);
  and g28 (n_185, in_0[6], in_0[7]);
  and g29 (n_69, in_1[0], in_1[1]);
  and g30 (n_71, in_1[0], in_1[2]);
  and g31 (n_73, in_1[1], in_1[2]);
  and g32 (n_72, in_1[0], in_1[3]);
  and g33 (n_81, in_1[1], in_1[3]);
  and g34 (n_89, in_1[2], in_1[3]);
  and g35 (n_80, in_1[0], in_1[4]);
  and g36 (n_91, in_1[1], in_1[4]);
  and g37 (n_100, in_1[2], in_1[4]);
  and g38 (n_66, in_1[3], in_1[4]);
  and g39 (n_88, in_1[0], in_1[5]);
  and g40 (n_49, in_1[1], in_1[5]);
  and g41 (n_111, in_1[2], in_1[5]);
  and g42 (n_126, in_1[3], in_1[5]);
  and g43 (n_144, in_1[4], in_1[5]);
  and g44 (n_51, in_1[0], in_1[6]);
  and g45 (n_112, in_1[1], in_1[6]);
  and g46 (n_127, in_1[2], in_1[6]);
  and g47 (n_146, in_1[3], in_1[6]);
  and g48 (n_160, in_1[4], in_1[6]);
  and g49 (n_169, in_1[5], in_1[6]);
  and g50 (n_114, in_1[0], in_1[7]);
  and g51 (n_129, in_1[1], in_1[7]);
  and g52 (n_143, in_1[2], in_1[7]);
  and g53 (n_159, in_1[3], in_1[7]);
  and g54 (n_172, in_1[4], in_1[7]);
  and g55 (n_180, in_1[5], in_1[7]);
  and g56 (n_186, in_1[6], in_1[7]);
  xor g106 (n_189, in_0[1], in_1[1]);
  xor g107 (n_65, n_189, n_69);
  nand g108 (n_190, in_0[1], in_1[1]);
  nand g109 (n_191, n_69, in_1[1]);
  nand g110 (n_192, in_0[1], n_69);
  nand g111 (n_64, n_190, n_191, n_192);
  xor g112 (n_47, n_70, n_71);
  and g113 (n_77, n_70, n_71);
  xor g114 (n_76, in_0[2], in_1[2]);
  and g115 (n_82, in_0[2], in_1[2]);
  xor g116 (n_193, n_72, n_73);
  xor g117 (n_46, n_193, n_74);
  nand g118 (n_194, n_72, n_73);
  nand g119 (n_195, n_74, n_73);
  nand g120 (n_196, n_72, n_74);
  nand g121 (n_84, n_194, n_195, n_196);
  xor g122 (n_197, n_75, n_76);
  xor g123 (n_63, n_197, n_77);
  nand g124 (n_198, n_75, n_76);
  nand g125 (n_199, n_77, n_76);
  nand g126 (n_200, n_75, n_77);
  nand g127 (n_45, n_198, n_199, n_200);
  xor g128 (n_83, n_78, n_79);
  and g129 (n_93, n_78, n_79);
  xor g130 (n_201, n_80, n_81);
  xor g131 (n_85, n_201, n_82);
  nand g132 (n_202, n_80, n_81);
  nand g133 (n_203, n_82, n_81);
  nand g134 (n_204, n_80, n_82);
  nand g135 (n_95, n_202, n_203, n_204);
  xor g136 (n_205, n_83, n_84);
  xor g137 (n_62, n_205, n_85);
  nand g138 (n_206, n_83, n_84);
  nand g139 (n_207, n_85, n_84);
  nand g140 (n_208, n_83, n_85);
  nand g141 (n_44, n_206, n_207, n_208);
  xor g142 (n_92, in_0[3], in_1[3]);
  and g143 (n_101, in_0[3], in_1[3]);
  xor g144 (n_209, n_86, n_87);
  xor g145 (n_96, n_209, n_88);
  nand g146 (n_210, n_86, n_87);
  nand g147 (n_211, n_88, n_87);
  nand g148 (n_212, n_86, n_88);
  nand g149 (n_103, n_210, n_211, n_212);
  xor g150 (n_213, n_89, n_90);
  xor g151 (n_94, n_213, n_91);
  nand g152 (n_214, n_89, n_90);
  nand g153 (n_215, n_91, n_90);
  nand g154 (n_216, n_89, n_91);
  nand g155 (n_104, n_214, n_215, n_216);
  xor g156 (n_217, n_92, n_93);
  xor g157 (n_97, n_217, n_94);
  nand g158 (n_218, n_92, n_93);
  nand g159 (n_219, n_94, n_93);
  nand g160 (n_220, n_92, n_94);
  nand g161 (n_108, n_218, n_219, n_220);
  xor g162 (n_221, n_95, n_96);
  xor g163 (n_61, n_221, n_97);
  nand g164 (n_222, n_95, n_96);
  nand g165 (n_223, n_97, n_96);
  nand g166 (n_224, n_95, n_97);
  nand g167 (n_43, n_222, n_223, n_224);
  xor g168 (n_102, n_98, n_99);
  and g169 (n_115, n_98, n_99);
  xor g170 (n_225, n_100, n_49);
  xor g171 (n_105, n_225, n_50);
  nand g172 (n_226, n_100, n_49);
  nand g173 (n_227, n_50, n_49);
  nand g174 (n_228, n_100, n_50);
  nand g175 (n_116, n_226, n_227, n_228);
  xor g176 (n_229, n_51, n_101);
  xor g177 (n_106, n_229, n_102);
  nand g178 (n_230, n_51, n_101);
  nand g179 (n_231, n_102, n_101);
  nand g180 (n_232, n_51, n_102);
  nand g181 (n_120, n_230, n_231, n_232);
  xor g182 (n_233, n_103, n_104);
  xor g183 (n_107, n_233, n_105);
  nand g184 (n_234, n_103, n_104);
  nand g185 (n_235, n_105, n_104);
  nand g186 (n_236, n_103, n_105);
  nand g187 (n_121, n_234, n_235, n_236);
  xor g188 (n_237, n_106, n_107);
  xor g189 (n_60, n_237, n_108);
  nand g190 (n_238, n_106, n_107);
  nand g191 (n_239, n_108, n_107);
  nand g192 (n_240, n_106, n_108);
  nand g193 (n_42, n_238, n_239, n_240);
  xor g194 (n_68, in_0[4], in_1[4]);
  and g195 (n_130, in_0[4], in_1[4]);
  xor g196 (n_241, n_109, n_110);
  xor g197 (n_117, n_241, n_111);
  nand g198 (n_242, n_109, n_110);
  nand g199 (n_243, n_111, n_110);
  nand g200 (n_244, n_109, n_111);
  nand g201 (n_133, n_242, n_243, n_244);
  xor g202 (n_245, n_112, n_113);
  xor g203 (n_119, n_245, n_114);
  nand g204 (n_246, n_112, n_113);
  nand g205 (n_247, n_114, n_113);
  nand g206 (n_248, n_112, n_114);
  nand g207 (n_132, n_246, n_247, n_248);
  xor g208 (n_249, n_66, n_67);
  xor g209 (n_118, n_249, n_68);
  nand g210 (n_250, n_66, n_67);
  nand g211 (n_251, n_68, n_67);
  nand g212 (n_252, n_66, n_68);
  nand g213 (n_134, n_250, n_251, n_252);
  xor g214 (n_253, n_115, n_116);
  xor g215 (n_122, n_253, n_117);
  nand g216 (n_254, n_115, n_116);
  nand g217 (n_255, n_117, n_116);
  nand g218 (n_256, n_115, n_117);
  nand g219 (n_138, n_254, n_255, n_256);
  xor g220 (n_257, n_118, n_119);
  xor g221 (n_123, n_257, n_120);
  nand g222 (n_258, n_118, n_119);
  nand g223 (n_259, n_120, n_119);
  nand g224 (n_260, n_118, n_120);
  nand g225 (n_139, n_258, n_259, n_260);
  xor g226 (n_261, n_121, n_122);
  xor g227 (n_59, n_261, n_123);
  nand g228 (n_262, n_121, n_122);
  nand g229 (n_263, n_123, n_122);
  nand g230 (n_264, n_121, n_123);
  nand g231 (n_41, n_262, n_263, n_264);
  xor g232 (n_131, n_124, n_125);
  and g233 (n_147, n_124, n_125);
  xor g234 (n_265, n_126, n_127);
  xor g235 (n_135, n_265, n_128);
  nand g236 (n_266, n_126, n_127);
  nand g237 (n_267, n_128, n_127);
  nand g238 (n_268, n_126, n_128);
  nand g239 (n_148, n_266, n_267, n_268);
  xor g240 (n_269, n_129, n_130);
  xor g241 (n_136, n_269, n_131);
  nand g242 (n_270, n_129, n_130);
  nand g243 (n_271, n_131, n_130);
  nand g244 (n_272, n_129, n_131);
  nand g245 (n_151, n_270, n_271, n_272);
  xor g246 (n_273, n_132, n_133);
  xor g247 (n_137, n_273, n_134);
  nand g248 (n_274, n_132, n_133);
  nand g249 (n_275, n_134, n_133);
  nand g250 (n_276, n_132, n_134);
  nand g251 (n_154, n_274, n_275, n_276);
  xor g252 (n_277, n_135, n_136);
  xor g253 (n_140, n_277, n_137);
  nand g254 (n_278, n_135, n_136);
  nand g255 (n_279, n_137, n_136);
  nand g256 (n_280, n_135, n_137);
  nand g257 (n_156, n_278, n_279, n_280);
  xor g258 (n_281, n_138, n_139);
  xor g259 (n_58, n_281, n_140);
  nand g260 (n_282, n_138, n_139);
  nand g261 (n_283, n_140, n_139);
  nand g262 (n_284, n_138, n_140);
  nand g263 (n_40, n_282, n_283, n_284);
  xor g264 (n_285, in_0[5], in_1[5]);
  xor g265 (n_149, n_285, n_141);
  nand g266 (n_286, in_0[5], in_1[5]);
  nand g267 (n_287, n_141, in_1[5]);
  nand g268 (n_288, in_0[5], n_141);
  nand g269 (n_161, n_286, n_287, n_288);
  xor g270 (n_289, n_142, n_143);
  xor g271 (n_150, n_289, n_144);
  nand g272 (n_290, n_142, n_143);
  nand g273 (n_291, n_144, n_143);
  nand g274 (n_292, n_142, n_144);
  nand g275 (n_162, n_290, n_291, n_292);
  xor g276 (n_293, n_145, n_146);
  xor g277 (n_152, n_293, n_147);
  nand g278 (n_294, n_145, n_146);
  nand g279 (n_295, n_147, n_146);
  nand g280 (n_296, n_145, n_147);
  nand g281 (n_164, n_294, n_295, n_296);
  xor g282 (n_297, n_148, n_149);
  xor g283 (n_153, n_297, n_150);
  nand g284 (n_298, n_148, n_149);
  nand g285 (n_299, n_150, n_149);
  nand g286 (n_300, n_148, n_150);
  nand g287 (n_165, n_298, n_299, n_300);
  xor g288 (n_301, n_151, n_152);
  xor g289 (n_155, n_301, n_153);
  nand g290 (n_302, n_151, n_152);
  nand g291 (n_303, n_153, n_152);
  nand g292 (n_304, n_151, n_153);
  nand g293 (n_168, n_302, n_303, n_304);
  xor g294 (n_305, n_154, n_155);
  xor g295 (n_57, n_305, n_156);
  nand g296 (n_306, n_154, n_155);
  nand g297 (n_307, n_156, n_155);
  nand g298 (n_308, n_154, n_156);
  nand g299 (n_39, n_306, n_307, n_308);
  xor g300 (n_309, n_157, n_158);
  xor g301 (n_163, n_309, n_159);
  nand g302 (n_310, n_157, n_158);
  nand g303 (n_311, n_159, n_158);
  nand g304 (n_312, n_157, n_159);
  nand g305 (n_174, n_310, n_311, n_312);
  xor g306 (n_313, n_160, n_161);
  xor g307 (n_166, n_313, n_162);
  nand g308 (n_314, n_160, n_161);
  nand g309 (n_315, n_162, n_161);
  nand g310 (n_316, n_160, n_162);
  nand g311 (n_176, n_314, n_315, n_316);
  xor g312 (n_317, n_163, n_164);
  xor g313 (n_167, n_317, n_165);
  nand g314 (n_318, n_163, n_164);
  nand g315 (n_319, n_165, n_164);
  nand g316 (n_320, n_163, n_165);
  nand g317 (n_178, n_318, n_319, n_320);
  xor g318 (n_321, n_166, n_167);
  xor g319 (n_56, n_321, n_168);
  nand g320 (n_322, n_166, n_167);
  nand g321 (n_323, n_168, n_167);
  nand g322 (n_324, n_166, n_168);
  nand g323 (n_38, n_322, n_323, n_324);
  xor g324 (n_325, in_0[6], in_1[6]);
  xor g325 (n_173, n_325, n_169);
  nand g326 (n_326, in_0[6], in_1[6]);
  nand g327 (n_327, n_169, in_1[6]);
  nand g328 (n_328, in_0[6], n_169);
  nand g329 (n_182, n_326, n_327, n_328);
  xor g330 (n_329, n_170, n_171);
  xor g331 (n_175, n_329, n_172);
  nand g332 (n_330, n_170, n_171);
  nand g333 (n_331, n_172, n_171);
  nand g334 (n_332, n_170, n_172);
  nand g335 (n_181, n_330, n_331, n_332);
  xor g336 (n_333, n_173, n_174);
  xor g337 (n_177, n_333, n_175);
  nand g338 (n_334, n_173, n_174);
  nand g339 (n_335, n_175, n_174);
  nand g340 (n_336, n_173, n_175);
  nand g341 (n_184, n_334, n_335, n_336);
  xor g342 (n_337, n_176, n_177);
  xor g343 (n_55, n_337, n_178);
  nand g344 (n_338, n_176, n_177);
  nand g345 (n_339, n_178, n_177);
  nand g346 (n_340, n_176, n_178);
  nand g347 (n_54, n_338, n_339, n_340);
  xor g348 (n_341, n_179, n_180);
  xor g349 (n_183, n_341, n_181);
  nand g350 (n_342, n_179, n_180);
  nand g351 (n_343, n_181, n_180);
  nand g352 (n_344, n_179, n_181);
  nand g353 (n_188, n_342, n_343, n_344);
  xor g354 (n_345, n_182, n_183);
  xor g355 (n_37, n_345, n_184);
  nand g356 (n_346, n_182, n_183);
  nand g357 (n_347, n_184, n_183);
  nand g358 (n_348, n_182, n_184);
  nand g359 (n_53, n_346, n_347, n_348);
  xor g360 (n_349, in_0[7], in_1[7]);
  xor g361 (n_187, n_349, n_185);
  nand g362 (n_350, in_0[7], in_1[7]);
  nand g363 (n_351, n_185, in_1[7]);
  nand g364 (n_352, in_0[7], n_185);
  nand g365 (n_35, n_350, n_351, n_352);
  xor g366 (n_353, n_186, n_187);
  xor g367 (n_36, n_353, n_188);
  nand g368 (n_354, n_186, n_187);
  nand g369 (n_355, n_188, n_187);
  nand g370 (n_356, n_186, n_188);
  nand g371 (n_52, n_354, n_355, n_356);
  nand g374 (n_358, in_1[0], in_0[0]);
  nor g379 (n_370, n_48, n_65);
  nand g380 (n_365, n_48, n_65);
  nor g381 (n_366, n_47, n_64);
  nand g382 (n_367, n_47, n_64);
  nor g383 (n_376, n_46, n_63);
  nand g384 (n_371, n_46, n_63);
  nor g385 (n_372, n_45, n_62);
  nand g386 (n_373, n_45, n_62);
  nor g387 (n_382, n_44, n_61);
  nand g388 (n_377, n_44, n_61);
  nor g389 (n_378, n_43, n_60);
  nand g390 (n_379, n_43, n_60);
  nor g391 (n_388, n_42, n_59);
  nand g392 (n_383, n_42, n_59);
  nor g393 (n_384, n_41, n_58);
  nand g394 (n_385, n_41, n_58);
  nor g395 (n_394, n_40, n_57);
  nand g396 (n_389, n_40, n_57);
  nor g397 (n_390, n_39, n_56);
  nand g398 (n_391, n_39, n_56);
  nor g399 (n_400, n_38, n_55);
  nand g400 (n_395, n_38, n_55);
  nor g401 (n_396, n_37, n_54);
  nand g402 (n_397, n_37, n_54);
  nor g403 (n_406, n_36, n_53);
  nand g404 (n_401, n_36, n_53);
  nor g405 (n_402, n_35, n_52);
  nand g406 (n_403, n_35, n_52);
  nor g412 (n_368, n_365, n_366);
  nor g416 (n_374, n_371, n_372);
  nor g419 (n_416, n_376, n_372);
  nor g420 (n_380, n_377, n_378);
  nor g423 (n_418, n_382, n_378);
  nor g424 (n_386, n_383, n_384);
  nor g427 (n_426, n_388, n_384);
  nor g57 (n_392, n_389, n_390);
  nor g60 (n_428, n_394, n_390);
  nor g61 (n_398, n_395, n_396);
  nor g64 (n_436, n_400, n_396);
  nor g65 (n_404, n_401, n_402);
  nor g68 (n_438, n_406, n_402);
  nor g74 (n_414, n_382, n_413);
  nand g83 (n_451, n_416, n_418);
  nor g84 (n_424, n_394, n_423);
  nand g93 (n_458, n_426, n_428);
  nor g94 (n_434, n_406, n_433);
  nand g103 (n_466, n_436, n_438);
  nand g428 (n_503, n_371, n_543);
  nand g430 (n_505, n_413, n_544);
  nand g433 (n_508, n_550, n_551);
  nand g436 (n_470, n_561, n_562);
  nor g437 (n_456, n_400, n_455);
  nor g440 (n_480, n_400, n_458);
  nor g446 (n_464, n_462, n_455);
  nor g449 (n_486, n_458, n_462);
  nor g450 (n_468, n_466, n_455);
  nor g453 (n_489, n_458, n_466);
  nand g456 (n_512, n_383, n_572);
  nand g457 (n_473, n_426, n_470);
  nand g458 (n_514, n_423, n_473);
  nand g461 (n_517, n_566, n_573);
  nand g464 (n_520, n_455, n_574);
  nand g465 (n_482, n_480, n_470);
  nand g466 (n_523, n_576, n_482);
  nand g467 (n_485, n_569, n_470);
  nand g468 (n_525, n_577, n_485);
  nand g469 (n_488, n_486, n_470);
  nand g470 (n_528, n_578, n_488);
  nand g471 (n_491, n_489, n_470);
  nand g472 (out_0[16], n_579, n_491);
  xnor g485 (out_0[5], n_503, n_546);
  xnor g487 (out_0[6], n_505, n_547);
  xnor g490 (out_0[7], n_508, n_552);
  xnor g492 (out_0[8], n_470, n_553);
  xnor g495 (out_0[9], n_512, n_558);
  xnor g497 (out_0[10], n_514, n_559);
  xnor g500 (out_0[11], n_517, n_563);
  xnor g503 (out_0[12], n_520, n_564);
  xnor g506 (out_0[13], n_523, n_565);
  xnor g508 (out_0[14], n_525, n_554);
  xnor g511 (out_0[15], n_528, n_555);
  xor g514 (out_0[0], in_0[0], in_1[0]);
  not g515 (out_0[1], n_358);
  or g516 (n_535, wc, n_370);
  not gc (wc, n_365);
  and g517 (n_536, wc0, n_367);
  not gc0 (wc0, n_368);
  not g519 (out_0[2], n_535);
  or g520 (n_539, wc1, n_366);
  not gc1 (wc1, n_367);
  or g521 (n_540, wc2, n_376);
  not gc2 (wc2, n_371);
  xor g523 (out_0[3], n_365, n_539);
  and g524 (n_413, wc3, n_373);
  not gc3 (wc3, n_374);
  or g525 (n_542, wc4, n_382);
  not gc4 (wc4, n_416);
  or g526 (n_543, n_376, n_536);
  or g527 (n_544, n_536, wc5);
  not gc5 (wc5, n_416);
  xor g528 (out_0[4], n_536, n_540);
  or g529 (n_546, wc6, n_372);
  not gc6 (wc6, n_373);
  or g530 (n_547, wc7, n_382);
  not gc7 (wc7, n_377);
  and g531 (n_548, wc8, n_379);
  not gc8 (wc8, n_380);
  and g532 (n_549, wc9, n_403);
  not gc9 (wc9, n_404);
  and g533 (n_550, wc10, n_377);
  not gc10 (wc10, n_414);
  or g534 (n_551, n_536, n_542);
  or g535 (n_552, wc11, n_378);
  not gc11 (wc11, n_379);
  or g536 (n_553, wc12, n_388);
  not gc12 (wc12, n_383);
  or g537 (n_554, wc13, n_406);
  not gc13 (wc13, n_401);
  or g538 (n_555, wc14, n_402);
  not gc14 (wc14, n_403);
  and g539 (n_423, wc15, n_385);
  not gc15 (wc15, n_386);
  and g540 (n_556, wc16, n_418);
  not gc16 (wc16, n_413);
  or g541 (n_557, wc17, n_394);
  not gc17 (wc17, n_426);
  or g542 (n_558, wc18, n_384);
  not gc18 (wc18, n_385);
  or g543 (n_559, wc19, n_394);
  not gc19 (wc19, n_389);
  and g544 (n_560, wc20, n_391);
  not gc20 (wc20, n_392);
  and g545 (n_433, wc21, n_397);
  not gc21 (wc21, n_398);
  and g546 (n_561, wc22, n_548);
  not gc22 (wc22, n_556);
  or g547 (n_462, wc23, n_406);
  not gc23 (wc23, n_436);
  or g548 (n_562, n_451, n_536);
  or g549 (n_563, wc24, n_390);
  not gc24 (wc24, n_391);
  or g550 (n_564, wc25, n_400);
  not gc25 (wc25, n_395);
  or g551 (n_565, wc26, n_396);
  not gc26 (wc26, n_397);
  and g552 (n_566, wc27, n_389);
  not gc27 (wc27, n_424);
  and g553 (n_567, wc28, n_428);
  not gc28 (wc28, n_423);
  and g554 (n_568, wc29, n_438);
  not gc29 (wc29, n_433);
  and g555 (n_569, wc30, n_436);
  not gc30 (wc30, n_458);
  and g556 (n_455, wc31, n_560);
  not gc31 (wc31, n_567);
  and g557 (n_570, wc32, n_401);
  not gc32 (wc32, n_434);
  and g558 (n_571, wc33, n_549);
  not gc33 (wc33, n_568);
  or g559 (n_572, wc34, n_388);
  not gc34 (wc34, n_470);
  or g560 (n_573, n_557, wc35);
  not gc35 (wc35, n_470);
  or g561 (n_574, wc36, n_458);
  not gc36 (wc36, n_470);
  and g562 (n_575, wc37, n_436);
  not gc37 (wc37, n_455);
  and g563 (n_576, wc38, n_395);
  not gc38 (wc38, n_456);
  and g564 (n_577, wc39, n_433);
  not gc39 (wc39, n_575);
  and g565 (n_578, n_570, wc40);
  not gc40 (wc40, n_464);
  and g566 (n_579, n_571, wc41);
  not gc41 (wc41, n_468);
endmodule

module csa_tree_distance3_add1031_group_333_GENERIC(in_0, in_1, out_0);
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  csa_tree_distance3_add1031_group_333_GENERIC_REAL g1(.in_0 (in_0),
       .in_1 (in_1), .out_0 (out_0));
endmodule

module csa_tree_distance4_add1030_group_335_GENERIC_REAL(in_0, in_1,
     out_0);
// synthesis_equation "assign out_0 = ( ( in_0 * in_0 )  + ( in_1 * in_1 )  )  ;"
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_358, n_365, n_366, n_367, n_368, n_370;
  wire n_371, n_372, n_373, n_374, n_376, n_377, n_378, n_379;
  wire n_380, n_382, n_383, n_384, n_385, n_386, n_388, n_389;
  wire n_390, n_391, n_392, n_394, n_395, n_396, n_397, n_398;
  wire n_400, n_401, n_402, n_403, n_404, n_406, n_413, n_414;
  wire n_416, n_418, n_423, n_424, n_426, n_428, n_433, n_434;
  wire n_436, n_438, n_451, n_455, n_456, n_458, n_462, n_464;
  wire n_466, n_468, n_470, n_473, n_480, n_482, n_485, n_486;
  wire n_488, n_489, n_491, n_503, n_505, n_508, n_512, n_514;
  wire n_517, n_520, n_523, n_525, n_528, n_535, n_536, n_539;
  wire n_540, n_542, n_543, n_544, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579;
  and g1 (n_48, in_0[0], in_0[1]);
  and g2 (n_70, in_0[0], in_0[2]);
  and g3 (n_74, in_0[1], in_0[2]);
  and g4 (n_75, in_0[0], in_0[3]);
  and g5 (n_78, in_0[1], in_0[3]);
  and g6 (n_86, in_0[2], in_0[3]);
  and g7 (n_79, in_0[0], in_0[4]);
  and g8 (n_90, in_0[1], in_0[4]);
  and g9 (n_98, in_0[2], in_0[4]);
  and g10 (n_109, in_0[3], in_0[4]);
  and g11 (n_87, in_0[0], in_0[5]);
  and g12 (n_99, in_0[1], in_0[5]);
  and g13 (n_67, in_0[2], in_0[5]);
  and g14 (n_124, in_0[3], in_0[5]);
  and g15 (n_141, in_0[4], in_0[5]);
  and g16 (n_50, in_0[0], in_0[6]);
  and g17 (n_110, in_0[1], in_0[6]);
  and g18 (n_125, in_0[2], in_0[6]);
  and g19 (n_145, in_0[3], in_0[6]);
  and g20 (n_157, in_0[4], in_0[6]);
  and g21 (n_170, in_0[5], in_0[6]);
  and g22 (n_113, in_0[0], in_0[7]);
  and g23 (n_128, in_0[1], in_0[7]);
  and g24 (n_142, in_0[2], in_0[7]);
  and g25 (n_158, in_0[3], in_0[7]);
  and g26 (n_171, in_0[4], in_0[7]);
  and g27 (n_179, in_0[5], in_0[7]);
  and g28 (n_185, in_0[6], in_0[7]);
  and g29 (n_69, in_1[0], in_1[1]);
  and g30 (n_71, in_1[0], in_1[2]);
  and g31 (n_73, in_1[1], in_1[2]);
  and g32 (n_72, in_1[0], in_1[3]);
  and g33 (n_81, in_1[1], in_1[3]);
  and g34 (n_89, in_1[2], in_1[3]);
  and g35 (n_80, in_1[0], in_1[4]);
  and g36 (n_91, in_1[1], in_1[4]);
  and g37 (n_100, in_1[2], in_1[4]);
  and g38 (n_66, in_1[3], in_1[4]);
  and g39 (n_88, in_1[0], in_1[5]);
  and g40 (n_49, in_1[1], in_1[5]);
  and g41 (n_111, in_1[2], in_1[5]);
  and g42 (n_126, in_1[3], in_1[5]);
  and g43 (n_144, in_1[4], in_1[5]);
  and g44 (n_51, in_1[0], in_1[6]);
  and g45 (n_112, in_1[1], in_1[6]);
  and g46 (n_127, in_1[2], in_1[6]);
  and g47 (n_146, in_1[3], in_1[6]);
  and g48 (n_160, in_1[4], in_1[6]);
  and g49 (n_169, in_1[5], in_1[6]);
  and g50 (n_114, in_1[0], in_1[7]);
  and g51 (n_129, in_1[1], in_1[7]);
  and g52 (n_143, in_1[2], in_1[7]);
  and g53 (n_159, in_1[3], in_1[7]);
  and g54 (n_172, in_1[4], in_1[7]);
  and g55 (n_180, in_1[5], in_1[7]);
  and g56 (n_186, in_1[6], in_1[7]);
  xor g106 (n_189, in_0[1], in_1[1]);
  xor g107 (n_65, n_189, n_69);
  nand g108 (n_190, in_0[1], in_1[1]);
  nand g109 (n_191, n_69, in_1[1]);
  nand g110 (n_192, in_0[1], n_69);
  nand g111 (n_64, n_190, n_191, n_192);
  xor g112 (n_47, n_70, n_71);
  and g113 (n_77, n_70, n_71);
  xor g114 (n_76, in_0[2], in_1[2]);
  and g115 (n_82, in_0[2], in_1[2]);
  xor g116 (n_193, n_72, n_73);
  xor g117 (n_46, n_193, n_74);
  nand g118 (n_194, n_72, n_73);
  nand g119 (n_195, n_74, n_73);
  nand g120 (n_196, n_72, n_74);
  nand g121 (n_84, n_194, n_195, n_196);
  xor g122 (n_197, n_75, n_76);
  xor g123 (n_63, n_197, n_77);
  nand g124 (n_198, n_75, n_76);
  nand g125 (n_199, n_77, n_76);
  nand g126 (n_200, n_75, n_77);
  nand g127 (n_45, n_198, n_199, n_200);
  xor g128 (n_83, n_78, n_79);
  and g129 (n_93, n_78, n_79);
  xor g130 (n_201, n_80, n_81);
  xor g131 (n_85, n_201, n_82);
  nand g132 (n_202, n_80, n_81);
  nand g133 (n_203, n_82, n_81);
  nand g134 (n_204, n_80, n_82);
  nand g135 (n_95, n_202, n_203, n_204);
  xor g136 (n_205, n_83, n_84);
  xor g137 (n_62, n_205, n_85);
  nand g138 (n_206, n_83, n_84);
  nand g139 (n_207, n_85, n_84);
  nand g140 (n_208, n_83, n_85);
  nand g141 (n_44, n_206, n_207, n_208);
  xor g142 (n_92, in_0[3], in_1[3]);
  and g143 (n_101, in_0[3], in_1[3]);
  xor g144 (n_209, n_86, n_87);
  xor g145 (n_96, n_209, n_88);
  nand g146 (n_210, n_86, n_87);
  nand g147 (n_211, n_88, n_87);
  nand g148 (n_212, n_86, n_88);
  nand g149 (n_103, n_210, n_211, n_212);
  xor g150 (n_213, n_89, n_90);
  xor g151 (n_94, n_213, n_91);
  nand g152 (n_214, n_89, n_90);
  nand g153 (n_215, n_91, n_90);
  nand g154 (n_216, n_89, n_91);
  nand g155 (n_104, n_214, n_215, n_216);
  xor g156 (n_217, n_92, n_93);
  xor g157 (n_97, n_217, n_94);
  nand g158 (n_218, n_92, n_93);
  nand g159 (n_219, n_94, n_93);
  nand g160 (n_220, n_92, n_94);
  nand g161 (n_108, n_218, n_219, n_220);
  xor g162 (n_221, n_95, n_96);
  xor g163 (n_61, n_221, n_97);
  nand g164 (n_222, n_95, n_96);
  nand g165 (n_223, n_97, n_96);
  nand g166 (n_224, n_95, n_97);
  nand g167 (n_43, n_222, n_223, n_224);
  xor g168 (n_102, n_98, n_99);
  and g169 (n_115, n_98, n_99);
  xor g170 (n_225, n_100, n_49);
  xor g171 (n_105, n_225, n_50);
  nand g172 (n_226, n_100, n_49);
  nand g173 (n_227, n_50, n_49);
  nand g174 (n_228, n_100, n_50);
  nand g175 (n_116, n_226, n_227, n_228);
  xor g176 (n_229, n_51, n_101);
  xor g177 (n_106, n_229, n_102);
  nand g178 (n_230, n_51, n_101);
  nand g179 (n_231, n_102, n_101);
  nand g180 (n_232, n_51, n_102);
  nand g181 (n_120, n_230, n_231, n_232);
  xor g182 (n_233, n_103, n_104);
  xor g183 (n_107, n_233, n_105);
  nand g184 (n_234, n_103, n_104);
  nand g185 (n_235, n_105, n_104);
  nand g186 (n_236, n_103, n_105);
  nand g187 (n_121, n_234, n_235, n_236);
  xor g188 (n_237, n_106, n_107);
  xor g189 (n_60, n_237, n_108);
  nand g190 (n_238, n_106, n_107);
  nand g191 (n_239, n_108, n_107);
  nand g192 (n_240, n_106, n_108);
  nand g193 (n_42, n_238, n_239, n_240);
  xor g194 (n_68, in_0[4], in_1[4]);
  and g195 (n_130, in_0[4], in_1[4]);
  xor g196 (n_241, n_109, n_110);
  xor g197 (n_117, n_241, n_111);
  nand g198 (n_242, n_109, n_110);
  nand g199 (n_243, n_111, n_110);
  nand g200 (n_244, n_109, n_111);
  nand g201 (n_133, n_242, n_243, n_244);
  xor g202 (n_245, n_112, n_113);
  xor g203 (n_119, n_245, n_114);
  nand g204 (n_246, n_112, n_113);
  nand g205 (n_247, n_114, n_113);
  nand g206 (n_248, n_112, n_114);
  nand g207 (n_132, n_246, n_247, n_248);
  xor g208 (n_249, n_66, n_67);
  xor g209 (n_118, n_249, n_68);
  nand g210 (n_250, n_66, n_67);
  nand g211 (n_251, n_68, n_67);
  nand g212 (n_252, n_66, n_68);
  nand g213 (n_134, n_250, n_251, n_252);
  xor g214 (n_253, n_115, n_116);
  xor g215 (n_122, n_253, n_117);
  nand g216 (n_254, n_115, n_116);
  nand g217 (n_255, n_117, n_116);
  nand g218 (n_256, n_115, n_117);
  nand g219 (n_138, n_254, n_255, n_256);
  xor g220 (n_257, n_118, n_119);
  xor g221 (n_123, n_257, n_120);
  nand g222 (n_258, n_118, n_119);
  nand g223 (n_259, n_120, n_119);
  nand g224 (n_260, n_118, n_120);
  nand g225 (n_139, n_258, n_259, n_260);
  xor g226 (n_261, n_121, n_122);
  xor g227 (n_59, n_261, n_123);
  nand g228 (n_262, n_121, n_122);
  nand g229 (n_263, n_123, n_122);
  nand g230 (n_264, n_121, n_123);
  nand g231 (n_41, n_262, n_263, n_264);
  xor g232 (n_131, n_124, n_125);
  and g233 (n_147, n_124, n_125);
  xor g234 (n_265, n_126, n_127);
  xor g235 (n_135, n_265, n_128);
  nand g236 (n_266, n_126, n_127);
  nand g237 (n_267, n_128, n_127);
  nand g238 (n_268, n_126, n_128);
  nand g239 (n_148, n_266, n_267, n_268);
  xor g240 (n_269, n_129, n_130);
  xor g241 (n_136, n_269, n_131);
  nand g242 (n_270, n_129, n_130);
  nand g243 (n_271, n_131, n_130);
  nand g244 (n_272, n_129, n_131);
  nand g245 (n_151, n_270, n_271, n_272);
  xor g246 (n_273, n_132, n_133);
  xor g247 (n_137, n_273, n_134);
  nand g248 (n_274, n_132, n_133);
  nand g249 (n_275, n_134, n_133);
  nand g250 (n_276, n_132, n_134);
  nand g251 (n_154, n_274, n_275, n_276);
  xor g252 (n_277, n_135, n_136);
  xor g253 (n_140, n_277, n_137);
  nand g254 (n_278, n_135, n_136);
  nand g255 (n_279, n_137, n_136);
  nand g256 (n_280, n_135, n_137);
  nand g257 (n_156, n_278, n_279, n_280);
  xor g258 (n_281, n_138, n_139);
  xor g259 (n_58, n_281, n_140);
  nand g260 (n_282, n_138, n_139);
  nand g261 (n_283, n_140, n_139);
  nand g262 (n_284, n_138, n_140);
  nand g263 (n_40, n_282, n_283, n_284);
  xor g264 (n_285, in_0[5], in_1[5]);
  xor g265 (n_149, n_285, n_141);
  nand g266 (n_286, in_0[5], in_1[5]);
  nand g267 (n_287, n_141, in_1[5]);
  nand g268 (n_288, in_0[5], n_141);
  nand g269 (n_161, n_286, n_287, n_288);
  xor g270 (n_289, n_142, n_143);
  xor g271 (n_150, n_289, n_144);
  nand g272 (n_290, n_142, n_143);
  nand g273 (n_291, n_144, n_143);
  nand g274 (n_292, n_142, n_144);
  nand g275 (n_162, n_290, n_291, n_292);
  xor g276 (n_293, n_145, n_146);
  xor g277 (n_152, n_293, n_147);
  nand g278 (n_294, n_145, n_146);
  nand g279 (n_295, n_147, n_146);
  nand g280 (n_296, n_145, n_147);
  nand g281 (n_164, n_294, n_295, n_296);
  xor g282 (n_297, n_148, n_149);
  xor g283 (n_153, n_297, n_150);
  nand g284 (n_298, n_148, n_149);
  nand g285 (n_299, n_150, n_149);
  nand g286 (n_300, n_148, n_150);
  nand g287 (n_165, n_298, n_299, n_300);
  xor g288 (n_301, n_151, n_152);
  xor g289 (n_155, n_301, n_153);
  nand g290 (n_302, n_151, n_152);
  nand g291 (n_303, n_153, n_152);
  nand g292 (n_304, n_151, n_153);
  nand g293 (n_168, n_302, n_303, n_304);
  xor g294 (n_305, n_154, n_155);
  xor g295 (n_57, n_305, n_156);
  nand g296 (n_306, n_154, n_155);
  nand g297 (n_307, n_156, n_155);
  nand g298 (n_308, n_154, n_156);
  nand g299 (n_39, n_306, n_307, n_308);
  xor g300 (n_309, n_157, n_158);
  xor g301 (n_163, n_309, n_159);
  nand g302 (n_310, n_157, n_158);
  nand g303 (n_311, n_159, n_158);
  nand g304 (n_312, n_157, n_159);
  nand g305 (n_174, n_310, n_311, n_312);
  xor g306 (n_313, n_160, n_161);
  xor g307 (n_166, n_313, n_162);
  nand g308 (n_314, n_160, n_161);
  nand g309 (n_315, n_162, n_161);
  nand g310 (n_316, n_160, n_162);
  nand g311 (n_176, n_314, n_315, n_316);
  xor g312 (n_317, n_163, n_164);
  xor g313 (n_167, n_317, n_165);
  nand g314 (n_318, n_163, n_164);
  nand g315 (n_319, n_165, n_164);
  nand g316 (n_320, n_163, n_165);
  nand g317 (n_178, n_318, n_319, n_320);
  xor g318 (n_321, n_166, n_167);
  xor g319 (n_56, n_321, n_168);
  nand g320 (n_322, n_166, n_167);
  nand g321 (n_323, n_168, n_167);
  nand g322 (n_324, n_166, n_168);
  nand g323 (n_38, n_322, n_323, n_324);
  xor g324 (n_325, in_0[6], in_1[6]);
  xor g325 (n_173, n_325, n_169);
  nand g326 (n_326, in_0[6], in_1[6]);
  nand g327 (n_327, n_169, in_1[6]);
  nand g328 (n_328, in_0[6], n_169);
  nand g329 (n_182, n_326, n_327, n_328);
  xor g330 (n_329, n_170, n_171);
  xor g331 (n_175, n_329, n_172);
  nand g332 (n_330, n_170, n_171);
  nand g333 (n_331, n_172, n_171);
  nand g334 (n_332, n_170, n_172);
  nand g335 (n_181, n_330, n_331, n_332);
  xor g336 (n_333, n_173, n_174);
  xor g337 (n_177, n_333, n_175);
  nand g338 (n_334, n_173, n_174);
  nand g339 (n_335, n_175, n_174);
  nand g340 (n_336, n_173, n_175);
  nand g341 (n_184, n_334, n_335, n_336);
  xor g342 (n_337, n_176, n_177);
  xor g343 (n_55, n_337, n_178);
  nand g344 (n_338, n_176, n_177);
  nand g345 (n_339, n_178, n_177);
  nand g346 (n_340, n_176, n_178);
  nand g347 (n_54, n_338, n_339, n_340);
  xor g348 (n_341, n_179, n_180);
  xor g349 (n_183, n_341, n_181);
  nand g350 (n_342, n_179, n_180);
  nand g351 (n_343, n_181, n_180);
  nand g352 (n_344, n_179, n_181);
  nand g353 (n_188, n_342, n_343, n_344);
  xor g354 (n_345, n_182, n_183);
  xor g355 (n_37, n_345, n_184);
  nand g356 (n_346, n_182, n_183);
  nand g357 (n_347, n_184, n_183);
  nand g358 (n_348, n_182, n_184);
  nand g359 (n_53, n_346, n_347, n_348);
  xor g360 (n_349, in_0[7], in_1[7]);
  xor g361 (n_187, n_349, n_185);
  nand g362 (n_350, in_0[7], in_1[7]);
  nand g363 (n_351, n_185, in_1[7]);
  nand g364 (n_352, in_0[7], n_185);
  nand g365 (n_35, n_350, n_351, n_352);
  xor g366 (n_353, n_186, n_187);
  xor g367 (n_36, n_353, n_188);
  nand g368 (n_354, n_186, n_187);
  nand g369 (n_355, n_188, n_187);
  nand g370 (n_356, n_186, n_188);
  nand g371 (n_52, n_354, n_355, n_356);
  nand g374 (n_358, in_1[0], in_0[0]);
  nor g379 (n_370, n_48, n_65);
  nand g380 (n_365, n_48, n_65);
  nor g381 (n_366, n_47, n_64);
  nand g382 (n_367, n_47, n_64);
  nor g383 (n_376, n_46, n_63);
  nand g384 (n_371, n_46, n_63);
  nor g385 (n_372, n_45, n_62);
  nand g386 (n_373, n_45, n_62);
  nor g387 (n_382, n_44, n_61);
  nand g388 (n_377, n_44, n_61);
  nor g389 (n_378, n_43, n_60);
  nand g390 (n_379, n_43, n_60);
  nor g391 (n_388, n_42, n_59);
  nand g392 (n_383, n_42, n_59);
  nor g393 (n_384, n_41, n_58);
  nand g394 (n_385, n_41, n_58);
  nor g395 (n_394, n_40, n_57);
  nand g396 (n_389, n_40, n_57);
  nor g397 (n_390, n_39, n_56);
  nand g398 (n_391, n_39, n_56);
  nor g399 (n_400, n_38, n_55);
  nand g400 (n_395, n_38, n_55);
  nor g401 (n_396, n_37, n_54);
  nand g402 (n_397, n_37, n_54);
  nor g403 (n_406, n_36, n_53);
  nand g404 (n_401, n_36, n_53);
  nor g405 (n_402, n_35, n_52);
  nand g406 (n_403, n_35, n_52);
  nor g412 (n_368, n_365, n_366);
  nor g416 (n_374, n_371, n_372);
  nor g419 (n_416, n_376, n_372);
  nor g420 (n_380, n_377, n_378);
  nor g423 (n_418, n_382, n_378);
  nor g424 (n_386, n_383, n_384);
  nor g427 (n_426, n_388, n_384);
  nor g57 (n_392, n_389, n_390);
  nor g60 (n_428, n_394, n_390);
  nor g61 (n_398, n_395, n_396);
  nor g64 (n_436, n_400, n_396);
  nor g65 (n_404, n_401, n_402);
  nor g68 (n_438, n_406, n_402);
  nor g74 (n_414, n_382, n_413);
  nand g83 (n_451, n_416, n_418);
  nor g84 (n_424, n_394, n_423);
  nand g93 (n_458, n_426, n_428);
  nor g94 (n_434, n_406, n_433);
  nand g103 (n_466, n_436, n_438);
  nand g428 (n_503, n_371, n_543);
  nand g430 (n_505, n_413, n_544);
  nand g433 (n_508, n_550, n_551);
  nand g436 (n_470, n_561, n_562);
  nor g437 (n_456, n_400, n_455);
  nor g440 (n_480, n_400, n_458);
  nor g446 (n_464, n_462, n_455);
  nor g449 (n_486, n_458, n_462);
  nor g450 (n_468, n_466, n_455);
  nor g453 (n_489, n_458, n_466);
  nand g456 (n_512, n_383, n_572);
  nand g457 (n_473, n_426, n_470);
  nand g458 (n_514, n_423, n_473);
  nand g461 (n_517, n_566, n_573);
  nand g464 (n_520, n_455, n_574);
  nand g465 (n_482, n_480, n_470);
  nand g466 (n_523, n_576, n_482);
  nand g467 (n_485, n_569, n_470);
  nand g468 (n_525, n_577, n_485);
  nand g469 (n_488, n_486, n_470);
  nand g470 (n_528, n_578, n_488);
  nand g471 (n_491, n_489, n_470);
  nand g472 (out_0[16], n_579, n_491);
  xnor g485 (out_0[5], n_503, n_546);
  xnor g487 (out_0[6], n_505, n_547);
  xnor g490 (out_0[7], n_508, n_552);
  xnor g492 (out_0[8], n_470, n_553);
  xnor g495 (out_0[9], n_512, n_558);
  xnor g497 (out_0[10], n_514, n_559);
  xnor g500 (out_0[11], n_517, n_563);
  xnor g503 (out_0[12], n_520, n_564);
  xnor g506 (out_0[13], n_523, n_565);
  xnor g508 (out_0[14], n_525, n_554);
  xnor g511 (out_0[15], n_528, n_555);
  xor g514 (out_0[0], in_0[0], in_1[0]);
  not g515 (out_0[1], n_358);
  or g516 (n_535, wc, n_370);
  not gc (wc, n_365);
  and g517 (n_536, wc0, n_367);
  not gc0 (wc0, n_368);
  not g519 (out_0[2], n_535);
  or g520 (n_539, wc1, n_366);
  not gc1 (wc1, n_367);
  or g521 (n_540, wc2, n_376);
  not gc2 (wc2, n_371);
  xor g523 (out_0[3], n_365, n_539);
  and g524 (n_413, wc3, n_373);
  not gc3 (wc3, n_374);
  or g525 (n_542, wc4, n_382);
  not gc4 (wc4, n_416);
  or g526 (n_543, n_376, n_536);
  or g527 (n_544, n_536, wc5);
  not gc5 (wc5, n_416);
  xor g528 (out_0[4], n_536, n_540);
  or g529 (n_546, wc6, n_372);
  not gc6 (wc6, n_373);
  or g530 (n_547, wc7, n_382);
  not gc7 (wc7, n_377);
  and g531 (n_548, wc8, n_379);
  not gc8 (wc8, n_380);
  and g532 (n_549, wc9, n_403);
  not gc9 (wc9, n_404);
  and g533 (n_550, wc10, n_377);
  not gc10 (wc10, n_414);
  or g534 (n_551, n_536, n_542);
  or g535 (n_552, wc11, n_378);
  not gc11 (wc11, n_379);
  or g536 (n_553, wc12, n_388);
  not gc12 (wc12, n_383);
  or g537 (n_554, wc13, n_406);
  not gc13 (wc13, n_401);
  or g538 (n_555, wc14, n_402);
  not gc14 (wc14, n_403);
  and g539 (n_423, wc15, n_385);
  not gc15 (wc15, n_386);
  and g540 (n_556, wc16, n_418);
  not gc16 (wc16, n_413);
  or g541 (n_557, wc17, n_394);
  not gc17 (wc17, n_426);
  or g542 (n_558, wc18, n_384);
  not gc18 (wc18, n_385);
  or g543 (n_559, wc19, n_394);
  not gc19 (wc19, n_389);
  and g544 (n_560, wc20, n_391);
  not gc20 (wc20, n_392);
  and g545 (n_433, wc21, n_397);
  not gc21 (wc21, n_398);
  and g546 (n_561, wc22, n_548);
  not gc22 (wc22, n_556);
  or g547 (n_462, wc23, n_406);
  not gc23 (wc23, n_436);
  or g548 (n_562, n_451, n_536);
  or g549 (n_563, wc24, n_390);
  not gc24 (wc24, n_391);
  or g550 (n_564, wc25, n_400);
  not gc25 (wc25, n_395);
  or g551 (n_565, wc26, n_396);
  not gc26 (wc26, n_397);
  and g552 (n_566, wc27, n_389);
  not gc27 (wc27, n_424);
  and g553 (n_567, wc28, n_428);
  not gc28 (wc28, n_423);
  and g554 (n_568, wc29, n_438);
  not gc29 (wc29, n_433);
  and g555 (n_569, wc30, n_436);
  not gc30 (wc30, n_458);
  and g556 (n_455, wc31, n_560);
  not gc31 (wc31, n_567);
  and g557 (n_570, wc32, n_401);
  not gc32 (wc32, n_434);
  and g558 (n_571, wc33, n_549);
  not gc33 (wc33, n_568);
  or g559 (n_572, wc34, n_388);
  not gc34 (wc34, n_470);
  or g560 (n_573, n_557, wc35);
  not gc35 (wc35, n_470);
  or g561 (n_574, wc36, n_458);
  not gc36 (wc36, n_470);
  and g562 (n_575, wc37, n_436);
  not gc37 (wc37, n_455);
  and g563 (n_576, wc38, n_395);
  not gc38 (wc38, n_456);
  and g564 (n_577, wc39, n_433);
  not gc39 (wc39, n_575);
  and g565 (n_578, n_570, wc40);
  not gc40 (wc40, n_464);
  and g566 (n_579, n_571, wc41);
  not gc41 (wc41, n_468);
endmodule

module csa_tree_distance4_add1030_group_335_GENERIC(in_0, in_1, out_0);
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  csa_tree_distance4_add1030_group_335_GENERIC_REAL g1(.in_0 (in_0),
       .in_1 (in_1), .out_0 (out_0));
endmodule

module csa_tree_distance5_add1029_group_337_GENERIC_REAL(in_0, in_1,
     out_0);
// synthesis_equation "assign out_0 = ( ( in_0 * in_0 )  + ( in_1 * in_1 )  )  ;"
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_358, n_365, n_366, n_367, n_368, n_370;
  wire n_371, n_372, n_373, n_374, n_376, n_377, n_378, n_379;
  wire n_380, n_382, n_383, n_384, n_385, n_386, n_388, n_389;
  wire n_390, n_391, n_392, n_394, n_395, n_396, n_397, n_398;
  wire n_400, n_401, n_402, n_403, n_404, n_406, n_413, n_414;
  wire n_416, n_418, n_423, n_424, n_426, n_428, n_433, n_434;
  wire n_436, n_438, n_451, n_455, n_456, n_458, n_462, n_464;
  wire n_466, n_468, n_470, n_473, n_480, n_482, n_485, n_486;
  wire n_488, n_489, n_491, n_503, n_505, n_508, n_512, n_514;
  wire n_517, n_520, n_523, n_525, n_528, n_535, n_536, n_539;
  wire n_540, n_542, n_543, n_544, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579;
  and g1 (n_48, in_0[0], in_0[1]);
  and g2 (n_70, in_0[0], in_0[2]);
  and g3 (n_74, in_0[1], in_0[2]);
  and g4 (n_75, in_0[0], in_0[3]);
  and g5 (n_78, in_0[1], in_0[3]);
  and g6 (n_86, in_0[2], in_0[3]);
  and g7 (n_79, in_0[0], in_0[4]);
  and g8 (n_90, in_0[1], in_0[4]);
  and g9 (n_98, in_0[2], in_0[4]);
  and g10 (n_109, in_0[3], in_0[4]);
  and g11 (n_87, in_0[0], in_0[5]);
  and g12 (n_99, in_0[1], in_0[5]);
  and g13 (n_67, in_0[2], in_0[5]);
  and g14 (n_124, in_0[3], in_0[5]);
  and g15 (n_141, in_0[4], in_0[5]);
  and g16 (n_50, in_0[0], in_0[6]);
  and g17 (n_110, in_0[1], in_0[6]);
  and g18 (n_125, in_0[2], in_0[6]);
  and g19 (n_145, in_0[3], in_0[6]);
  and g20 (n_157, in_0[4], in_0[6]);
  and g21 (n_170, in_0[5], in_0[6]);
  and g22 (n_113, in_0[0], in_0[7]);
  and g23 (n_128, in_0[1], in_0[7]);
  and g24 (n_142, in_0[2], in_0[7]);
  and g25 (n_158, in_0[3], in_0[7]);
  and g26 (n_171, in_0[4], in_0[7]);
  and g27 (n_179, in_0[5], in_0[7]);
  and g28 (n_185, in_0[6], in_0[7]);
  and g29 (n_69, in_1[0], in_1[1]);
  and g30 (n_71, in_1[0], in_1[2]);
  and g31 (n_73, in_1[1], in_1[2]);
  and g32 (n_72, in_1[0], in_1[3]);
  and g33 (n_81, in_1[1], in_1[3]);
  and g34 (n_89, in_1[2], in_1[3]);
  and g35 (n_80, in_1[0], in_1[4]);
  and g36 (n_91, in_1[1], in_1[4]);
  and g37 (n_100, in_1[2], in_1[4]);
  and g38 (n_66, in_1[3], in_1[4]);
  and g39 (n_88, in_1[0], in_1[5]);
  and g40 (n_49, in_1[1], in_1[5]);
  and g41 (n_111, in_1[2], in_1[5]);
  and g42 (n_126, in_1[3], in_1[5]);
  and g43 (n_144, in_1[4], in_1[5]);
  and g44 (n_51, in_1[0], in_1[6]);
  and g45 (n_112, in_1[1], in_1[6]);
  and g46 (n_127, in_1[2], in_1[6]);
  and g47 (n_146, in_1[3], in_1[6]);
  and g48 (n_160, in_1[4], in_1[6]);
  and g49 (n_169, in_1[5], in_1[6]);
  and g50 (n_114, in_1[0], in_1[7]);
  and g51 (n_129, in_1[1], in_1[7]);
  and g52 (n_143, in_1[2], in_1[7]);
  and g53 (n_159, in_1[3], in_1[7]);
  and g54 (n_172, in_1[4], in_1[7]);
  and g55 (n_180, in_1[5], in_1[7]);
  and g56 (n_186, in_1[6], in_1[7]);
  xor g106 (n_189, in_0[1], in_1[1]);
  xor g107 (n_65, n_189, n_69);
  nand g108 (n_190, in_0[1], in_1[1]);
  nand g109 (n_191, n_69, in_1[1]);
  nand g110 (n_192, in_0[1], n_69);
  nand g111 (n_64, n_190, n_191, n_192);
  xor g112 (n_47, n_70, n_71);
  and g113 (n_77, n_70, n_71);
  xor g114 (n_76, in_0[2], in_1[2]);
  and g115 (n_82, in_0[2], in_1[2]);
  xor g116 (n_193, n_72, n_73);
  xor g117 (n_46, n_193, n_74);
  nand g118 (n_194, n_72, n_73);
  nand g119 (n_195, n_74, n_73);
  nand g120 (n_196, n_72, n_74);
  nand g121 (n_84, n_194, n_195, n_196);
  xor g122 (n_197, n_75, n_76);
  xor g123 (n_63, n_197, n_77);
  nand g124 (n_198, n_75, n_76);
  nand g125 (n_199, n_77, n_76);
  nand g126 (n_200, n_75, n_77);
  nand g127 (n_45, n_198, n_199, n_200);
  xor g128 (n_83, n_78, n_79);
  and g129 (n_93, n_78, n_79);
  xor g130 (n_201, n_80, n_81);
  xor g131 (n_85, n_201, n_82);
  nand g132 (n_202, n_80, n_81);
  nand g133 (n_203, n_82, n_81);
  nand g134 (n_204, n_80, n_82);
  nand g135 (n_95, n_202, n_203, n_204);
  xor g136 (n_205, n_83, n_84);
  xor g137 (n_62, n_205, n_85);
  nand g138 (n_206, n_83, n_84);
  nand g139 (n_207, n_85, n_84);
  nand g140 (n_208, n_83, n_85);
  nand g141 (n_44, n_206, n_207, n_208);
  xor g142 (n_92, in_0[3], in_1[3]);
  and g143 (n_101, in_0[3], in_1[3]);
  xor g144 (n_209, n_86, n_87);
  xor g145 (n_96, n_209, n_88);
  nand g146 (n_210, n_86, n_87);
  nand g147 (n_211, n_88, n_87);
  nand g148 (n_212, n_86, n_88);
  nand g149 (n_103, n_210, n_211, n_212);
  xor g150 (n_213, n_89, n_90);
  xor g151 (n_94, n_213, n_91);
  nand g152 (n_214, n_89, n_90);
  nand g153 (n_215, n_91, n_90);
  nand g154 (n_216, n_89, n_91);
  nand g155 (n_104, n_214, n_215, n_216);
  xor g156 (n_217, n_92, n_93);
  xor g157 (n_97, n_217, n_94);
  nand g158 (n_218, n_92, n_93);
  nand g159 (n_219, n_94, n_93);
  nand g160 (n_220, n_92, n_94);
  nand g161 (n_108, n_218, n_219, n_220);
  xor g162 (n_221, n_95, n_96);
  xor g163 (n_61, n_221, n_97);
  nand g164 (n_222, n_95, n_96);
  nand g165 (n_223, n_97, n_96);
  nand g166 (n_224, n_95, n_97);
  nand g167 (n_43, n_222, n_223, n_224);
  xor g168 (n_102, n_98, n_99);
  and g169 (n_115, n_98, n_99);
  xor g170 (n_225, n_100, n_49);
  xor g171 (n_105, n_225, n_50);
  nand g172 (n_226, n_100, n_49);
  nand g173 (n_227, n_50, n_49);
  nand g174 (n_228, n_100, n_50);
  nand g175 (n_116, n_226, n_227, n_228);
  xor g176 (n_229, n_51, n_101);
  xor g177 (n_106, n_229, n_102);
  nand g178 (n_230, n_51, n_101);
  nand g179 (n_231, n_102, n_101);
  nand g180 (n_232, n_51, n_102);
  nand g181 (n_120, n_230, n_231, n_232);
  xor g182 (n_233, n_103, n_104);
  xor g183 (n_107, n_233, n_105);
  nand g184 (n_234, n_103, n_104);
  nand g185 (n_235, n_105, n_104);
  nand g186 (n_236, n_103, n_105);
  nand g187 (n_121, n_234, n_235, n_236);
  xor g188 (n_237, n_106, n_107);
  xor g189 (n_60, n_237, n_108);
  nand g190 (n_238, n_106, n_107);
  nand g191 (n_239, n_108, n_107);
  nand g192 (n_240, n_106, n_108);
  nand g193 (n_42, n_238, n_239, n_240);
  xor g194 (n_68, in_0[4], in_1[4]);
  and g195 (n_130, in_0[4], in_1[4]);
  xor g196 (n_241, n_109, n_110);
  xor g197 (n_117, n_241, n_111);
  nand g198 (n_242, n_109, n_110);
  nand g199 (n_243, n_111, n_110);
  nand g200 (n_244, n_109, n_111);
  nand g201 (n_133, n_242, n_243, n_244);
  xor g202 (n_245, n_112, n_113);
  xor g203 (n_119, n_245, n_114);
  nand g204 (n_246, n_112, n_113);
  nand g205 (n_247, n_114, n_113);
  nand g206 (n_248, n_112, n_114);
  nand g207 (n_132, n_246, n_247, n_248);
  xor g208 (n_249, n_66, n_67);
  xor g209 (n_118, n_249, n_68);
  nand g210 (n_250, n_66, n_67);
  nand g211 (n_251, n_68, n_67);
  nand g212 (n_252, n_66, n_68);
  nand g213 (n_134, n_250, n_251, n_252);
  xor g214 (n_253, n_115, n_116);
  xor g215 (n_122, n_253, n_117);
  nand g216 (n_254, n_115, n_116);
  nand g217 (n_255, n_117, n_116);
  nand g218 (n_256, n_115, n_117);
  nand g219 (n_138, n_254, n_255, n_256);
  xor g220 (n_257, n_118, n_119);
  xor g221 (n_123, n_257, n_120);
  nand g222 (n_258, n_118, n_119);
  nand g223 (n_259, n_120, n_119);
  nand g224 (n_260, n_118, n_120);
  nand g225 (n_139, n_258, n_259, n_260);
  xor g226 (n_261, n_121, n_122);
  xor g227 (n_59, n_261, n_123);
  nand g228 (n_262, n_121, n_122);
  nand g229 (n_263, n_123, n_122);
  nand g230 (n_264, n_121, n_123);
  nand g231 (n_41, n_262, n_263, n_264);
  xor g232 (n_131, n_124, n_125);
  and g233 (n_147, n_124, n_125);
  xor g234 (n_265, n_126, n_127);
  xor g235 (n_135, n_265, n_128);
  nand g236 (n_266, n_126, n_127);
  nand g237 (n_267, n_128, n_127);
  nand g238 (n_268, n_126, n_128);
  nand g239 (n_148, n_266, n_267, n_268);
  xor g240 (n_269, n_129, n_130);
  xor g241 (n_136, n_269, n_131);
  nand g242 (n_270, n_129, n_130);
  nand g243 (n_271, n_131, n_130);
  nand g244 (n_272, n_129, n_131);
  nand g245 (n_151, n_270, n_271, n_272);
  xor g246 (n_273, n_132, n_133);
  xor g247 (n_137, n_273, n_134);
  nand g248 (n_274, n_132, n_133);
  nand g249 (n_275, n_134, n_133);
  nand g250 (n_276, n_132, n_134);
  nand g251 (n_154, n_274, n_275, n_276);
  xor g252 (n_277, n_135, n_136);
  xor g253 (n_140, n_277, n_137);
  nand g254 (n_278, n_135, n_136);
  nand g255 (n_279, n_137, n_136);
  nand g256 (n_280, n_135, n_137);
  nand g257 (n_156, n_278, n_279, n_280);
  xor g258 (n_281, n_138, n_139);
  xor g259 (n_58, n_281, n_140);
  nand g260 (n_282, n_138, n_139);
  nand g261 (n_283, n_140, n_139);
  nand g262 (n_284, n_138, n_140);
  nand g263 (n_40, n_282, n_283, n_284);
  xor g264 (n_285, in_0[5], in_1[5]);
  xor g265 (n_149, n_285, n_141);
  nand g266 (n_286, in_0[5], in_1[5]);
  nand g267 (n_287, n_141, in_1[5]);
  nand g268 (n_288, in_0[5], n_141);
  nand g269 (n_161, n_286, n_287, n_288);
  xor g270 (n_289, n_142, n_143);
  xor g271 (n_150, n_289, n_144);
  nand g272 (n_290, n_142, n_143);
  nand g273 (n_291, n_144, n_143);
  nand g274 (n_292, n_142, n_144);
  nand g275 (n_162, n_290, n_291, n_292);
  xor g276 (n_293, n_145, n_146);
  xor g277 (n_152, n_293, n_147);
  nand g278 (n_294, n_145, n_146);
  nand g279 (n_295, n_147, n_146);
  nand g280 (n_296, n_145, n_147);
  nand g281 (n_164, n_294, n_295, n_296);
  xor g282 (n_297, n_148, n_149);
  xor g283 (n_153, n_297, n_150);
  nand g284 (n_298, n_148, n_149);
  nand g285 (n_299, n_150, n_149);
  nand g286 (n_300, n_148, n_150);
  nand g287 (n_165, n_298, n_299, n_300);
  xor g288 (n_301, n_151, n_152);
  xor g289 (n_155, n_301, n_153);
  nand g290 (n_302, n_151, n_152);
  nand g291 (n_303, n_153, n_152);
  nand g292 (n_304, n_151, n_153);
  nand g293 (n_168, n_302, n_303, n_304);
  xor g294 (n_305, n_154, n_155);
  xor g295 (n_57, n_305, n_156);
  nand g296 (n_306, n_154, n_155);
  nand g297 (n_307, n_156, n_155);
  nand g298 (n_308, n_154, n_156);
  nand g299 (n_39, n_306, n_307, n_308);
  xor g300 (n_309, n_157, n_158);
  xor g301 (n_163, n_309, n_159);
  nand g302 (n_310, n_157, n_158);
  nand g303 (n_311, n_159, n_158);
  nand g304 (n_312, n_157, n_159);
  nand g305 (n_174, n_310, n_311, n_312);
  xor g306 (n_313, n_160, n_161);
  xor g307 (n_166, n_313, n_162);
  nand g308 (n_314, n_160, n_161);
  nand g309 (n_315, n_162, n_161);
  nand g310 (n_316, n_160, n_162);
  nand g311 (n_176, n_314, n_315, n_316);
  xor g312 (n_317, n_163, n_164);
  xor g313 (n_167, n_317, n_165);
  nand g314 (n_318, n_163, n_164);
  nand g315 (n_319, n_165, n_164);
  nand g316 (n_320, n_163, n_165);
  nand g317 (n_178, n_318, n_319, n_320);
  xor g318 (n_321, n_166, n_167);
  xor g319 (n_56, n_321, n_168);
  nand g320 (n_322, n_166, n_167);
  nand g321 (n_323, n_168, n_167);
  nand g322 (n_324, n_166, n_168);
  nand g323 (n_38, n_322, n_323, n_324);
  xor g324 (n_325, in_0[6], in_1[6]);
  xor g325 (n_173, n_325, n_169);
  nand g326 (n_326, in_0[6], in_1[6]);
  nand g327 (n_327, n_169, in_1[6]);
  nand g328 (n_328, in_0[6], n_169);
  nand g329 (n_182, n_326, n_327, n_328);
  xor g330 (n_329, n_170, n_171);
  xor g331 (n_175, n_329, n_172);
  nand g332 (n_330, n_170, n_171);
  nand g333 (n_331, n_172, n_171);
  nand g334 (n_332, n_170, n_172);
  nand g335 (n_181, n_330, n_331, n_332);
  xor g336 (n_333, n_173, n_174);
  xor g337 (n_177, n_333, n_175);
  nand g338 (n_334, n_173, n_174);
  nand g339 (n_335, n_175, n_174);
  nand g340 (n_336, n_173, n_175);
  nand g341 (n_184, n_334, n_335, n_336);
  xor g342 (n_337, n_176, n_177);
  xor g343 (n_55, n_337, n_178);
  nand g344 (n_338, n_176, n_177);
  nand g345 (n_339, n_178, n_177);
  nand g346 (n_340, n_176, n_178);
  nand g347 (n_54, n_338, n_339, n_340);
  xor g348 (n_341, n_179, n_180);
  xor g349 (n_183, n_341, n_181);
  nand g350 (n_342, n_179, n_180);
  nand g351 (n_343, n_181, n_180);
  nand g352 (n_344, n_179, n_181);
  nand g353 (n_188, n_342, n_343, n_344);
  xor g354 (n_345, n_182, n_183);
  xor g355 (n_37, n_345, n_184);
  nand g356 (n_346, n_182, n_183);
  nand g357 (n_347, n_184, n_183);
  nand g358 (n_348, n_182, n_184);
  nand g359 (n_53, n_346, n_347, n_348);
  xor g360 (n_349, in_0[7], in_1[7]);
  xor g361 (n_187, n_349, n_185);
  nand g362 (n_350, in_0[7], in_1[7]);
  nand g363 (n_351, n_185, in_1[7]);
  nand g364 (n_352, in_0[7], n_185);
  nand g365 (n_35, n_350, n_351, n_352);
  xor g366 (n_353, n_186, n_187);
  xor g367 (n_36, n_353, n_188);
  nand g368 (n_354, n_186, n_187);
  nand g369 (n_355, n_188, n_187);
  nand g370 (n_356, n_186, n_188);
  nand g371 (n_52, n_354, n_355, n_356);
  nand g374 (n_358, in_1[0], in_0[0]);
  nor g379 (n_370, n_48, n_65);
  nand g380 (n_365, n_48, n_65);
  nor g381 (n_366, n_47, n_64);
  nand g382 (n_367, n_47, n_64);
  nor g383 (n_376, n_46, n_63);
  nand g384 (n_371, n_46, n_63);
  nor g385 (n_372, n_45, n_62);
  nand g386 (n_373, n_45, n_62);
  nor g387 (n_382, n_44, n_61);
  nand g388 (n_377, n_44, n_61);
  nor g389 (n_378, n_43, n_60);
  nand g390 (n_379, n_43, n_60);
  nor g391 (n_388, n_42, n_59);
  nand g392 (n_383, n_42, n_59);
  nor g393 (n_384, n_41, n_58);
  nand g394 (n_385, n_41, n_58);
  nor g395 (n_394, n_40, n_57);
  nand g396 (n_389, n_40, n_57);
  nor g397 (n_390, n_39, n_56);
  nand g398 (n_391, n_39, n_56);
  nor g399 (n_400, n_38, n_55);
  nand g400 (n_395, n_38, n_55);
  nor g401 (n_396, n_37, n_54);
  nand g402 (n_397, n_37, n_54);
  nor g403 (n_406, n_36, n_53);
  nand g404 (n_401, n_36, n_53);
  nor g405 (n_402, n_35, n_52);
  nand g406 (n_403, n_35, n_52);
  nor g412 (n_368, n_365, n_366);
  nor g416 (n_374, n_371, n_372);
  nor g419 (n_416, n_376, n_372);
  nor g420 (n_380, n_377, n_378);
  nor g423 (n_418, n_382, n_378);
  nor g424 (n_386, n_383, n_384);
  nor g427 (n_426, n_388, n_384);
  nor g57 (n_392, n_389, n_390);
  nor g60 (n_428, n_394, n_390);
  nor g61 (n_398, n_395, n_396);
  nor g64 (n_436, n_400, n_396);
  nor g65 (n_404, n_401, n_402);
  nor g68 (n_438, n_406, n_402);
  nor g74 (n_414, n_382, n_413);
  nand g83 (n_451, n_416, n_418);
  nor g84 (n_424, n_394, n_423);
  nand g93 (n_458, n_426, n_428);
  nor g94 (n_434, n_406, n_433);
  nand g103 (n_466, n_436, n_438);
  nand g428 (n_503, n_371, n_543);
  nand g430 (n_505, n_413, n_544);
  nand g433 (n_508, n_550, n_551);
  nand g436 (n_470, n_561, n_562);
  nor g437 (n_456, n_400, n_455);
  nor g440 (n_480, n_400, n_458);
  nor g446 (n_464, n_462, n_455);
  nor g449 (n_486, n_458, n_462);
  nor g450 (n_468, n_466, n_455);
  nor g453 (n_489, n_458, n_466);
  nand g456 (n_512, n_383, n_572);
  nand g457 (n_473, n_426, n_470);
  nand g458 (n_514, n_423, n_473);
  nand g461 (n_517, n_566, n_573);
  nand g464 (n_520, n_455, n_574);
  nand g465 (n_482, n_480, n_470);
  nand g466 (n_523, n_576, n_482);
  nand g467 (n_485, n_569, n_470);
  nand g468 (n_525, n_577, n_485);
  nand g469 (n_488, n_486, n_470);
  nand g470 (n_528, n_578, n_488);
  nand g471 (n_491, n_489, n_470);
  nand g472 (out_0[16], n_579, n_491);
  xnor g485 (out_0[5], n_503, n_546);
  xnor g487 (out_0[6], n_505, n_547);
  xnor g490 (out_0[7], n_508, n_552);
  xnor g492 (out_0[8], n_470, n_553);
  xnor g495 (out_0[9], n_512, n_558);
  xnor g497 (out_0[10], n_514, n_559);
  xnor g500 (out_0[11], n_517, n_563);
  xnor g503 (out_0[12], n_520, n_564);
  xnor g506 (out_0[13], n_523, n_565);
  xnor g508 (out_0[14], n_525, n_554);
  xnor g511 (out_0[15], n_528, n_555);
  xor g514 (out_0[0], in_0[0], in_1[0]);
  not g515 (out_0[1], n_358);
  or g516 (n_535, wc, n_370);
  not gc (wc, n_365);
  and g517 (n_536, wc0, n_367);
  not gc0 (wc0, n_368);
  not g519 (out_0[2], n_535);
  or g520 (n_539, wc1, n_366);
  not gc1 (wc1, n_367);
  or g521 (n_540, wc2, n_376);
  not gc2 (wc2, n_371);
  xor g523 (out_0[3], n_365, n_539);
  and g524 (n_413, wc3, n_373);
  not gc3 (wc3, n_374);
  or g525 (n_542, wc4, n_382);
  not gc4 (wc4, n_416);
  or g526 (n_543, n_376, n_536);
  or g527 (n_544, n_536, wc5);
  not gc5 (wc5, n_416);
  xor g528 (out_0[4], n_536, n_540);
  or g529 (n_546, wc6, n_372);
  not gc6 (wc6, n_373);
  or g530 (n_547, wc7, n_382);
  not gc7 (wc7, n_377);
  and g531 (n_548, wc8, n_379);
  not gc8 (wc8, n_380);
  and g532 (n_549, wc9, n_403);
  not gc9 (wc9, n_404);
  and g533 (n_550, wc10, n_377);
  not gc10 (wc10, n_414);
  or g534 (n_551, n_536, n_542);
  or g535 (n_552, wc11, n_378);
  not gc11 (wc11, n_379);
  or g536 (n_553, wc12, n_388);
  not gc12 (wc12, n_383);
  or g537 (n_554, wc13, n_406);
  not gc13 (wc13, n_401);
  or g538 (n_555, wc14, n_402);
  not gc14 (wc14, n_403);
  and g539 (n_423, wc15, n_385);
  not gc15 (wc15, n_386);
  and g540 (n_556, wc16, n_418);
  not gc16 (wc16, n_413);
  or g541 (n_557, wc17, n_394);
  not gc17 (wc17, n_426);
  or g542 (n_558, wc18, n_384);
  not gc18 (wc18, n_385);
  or g543 (n_559, wc19, n_394);
  not gc19 (wc19, n_389);
  and g544 (n_560, wc20, n_391);
  not gc20 (wc20, n_392);
  and g545 (n_433, wc21, n_397);
  not gc21 (wc21, n_398);
  and g546 (n_561, wc22, n_548);
  not gc22 (wc22, n_556);
  or g547 (n_462, wc23, n_406);
  not gc23 (wc23, n_436);
  or g548 (n_562, n_451, n_536);
  or g549 (n_563, wc24, n_390);
  not gc24 (wc24, n_391);
  or g550 (n_564, wc25, n_400);
  not gc25 (wc25, n_395);
  or g551 (n_565, wc26, n_396);
  not gc26 (wc26, n_397);
  and g552 (n_566, wc27, n_389);
  not gc27 (wc27, n_424);
  and g553 (n_567, wc28, n_428);
  not gc28 (wc28, n_423);
  and g554 (n_568, wc29, n_438);
  not gc29 (wc29, n_433);
  and g555 (n_569, wc30, n_436);
  not gc30 (wc30, n_458);
  and g556 (n_455, wc31, n_560);
  not gc31 (wc31, n_567);
  and g557 (n_570, wc32, n_401);
  not gc32 (wc32, n_434);
  and g558 (n_571, wc33, n_549);
  not gc33 (wc33, n_568);
  or g559 (n_572, wc34, n_388);
  not gc34 (wc34, n_470);
  or g560 (n_573, n_557, wc35);
  not gc35 (wc35, n_470);
  or g561 (n_574, wc36, n_458);
  not gc36 (wc36, n_470);
  and g562 (n_575, wc37, n_436);
  not gc37 (wc37, n_455);
  and g563 (n_576, wc38, n_395);
  not gc38 (wc38, n_456);
  and g564 (n_577, wc39, n_433);
  not gc39 (wc39, n_575);
  and g565 (n_578, n_570, wc40);
  not gc40 (wc40, n_464);
  and g566 (n_579, n_571, wc41);
  not gc41 (wc41, n_468);
endmodule

module csa_tree_distance5_add1029_group_337_GENERIC(in_0, in_1, out_0);
  input [7:0] in_0, in_1;
  output [16:0] out_0;
  wire [7:0] in_0, in_1;
  wire [16:0] out_0;
  csa_tree_distance5_add1029_group_337_GENERIC_REAL g1(.in_0 (in_0),
       .in_1 (in_1), .out_0 (out_0));
endmodule

module divide_unsigned_GENERIC_REAL(A, B, QUOTIENT);
// synthesis_equation "assign QUOTIENT = A / B;"
  input [14:0] A;
  input [6:0] B;
  output [14:0] QUOTIENT;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] QUOTIENT;
  wire n_39, n_40, n_42, n_43, n_44, n_45, n_46, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_56, n_57, n_59;
  wire n_60, n_63, n_64, n_65, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_80;
  wire n_81, n_82, n_85, n_86, n_87, n_88, n_89, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_110, n_111, n_112, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_147, n_150, n_151, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_165, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_192, n_195;
  wire n_196, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_210, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_237, n_240, n_241, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_286, n_302, n_305, n_308, n_310;
  wire n_311, n_312, n_313, n_316, n_317, n_318, n_319, n_322;
  wire n_325, n_327, n_329, n_331, n_332, n_335, n_336, n_342;
  wire n_346, n_348, n_349, n_358, n_360, n_377, n_379, n_381;
  wire n_382, n_383, n_384, n_387, n_388, n_408, n_411, n_413;
  wire n_414, n_415, n_416, n_419, n_420, n_431, n_448, n_450;
  wire n_451, n_452, n_453, n_456, n_457, n_458, n_460, n_468;
  wire n_487, n_489, n_491, n_493, n_494, n_495, n_496, n_498;
  wire n_499, n_500, n_501, n_502, n_505, n_507, n_510, n_512;
  wire n_522, n_535, n_536, n_539, n_541, n_542, n_543, n_544;
  wire n_546, n_547, n_548, n_549, n_550, n_553, n_555, n_558;
  wire n_563, n_570, n_576, n_594, n_596, n_597, n_598, n_599;
  wire n_601, n_602, n_603, n_604, n_605, n_608, n_610, n_613;
  wire n_618, n_625, n_633, n_650, n_652, n_654, n_656, n_657;
  wire n_658, n_659, n_661, n_662, n_663, n_664, n_665, n_667;
  wire n_668, n_671, n_673, n_674, n_675, n_676, n_677, n_679;
  wire n_681, n_684, n_692, n_696, n_698, n_709, n_710, n_713;
  wire n_715, n_716, n_717, n_718, n_720, n_721, n_722, n_723;
  wire n_724, n_726, n_727, n_728, n_729, n_730, n_733, n_735;
  wire n_736, n_739, n_741, n_744, n_747, n_752, n_754, n_759;
  wire n_763, n_765, n_780, n_782, n_783, n_784, n_785, n_787;
  wire n_788, n_789, n_790, n_791, n_793, n_794, n_795, n_796;
  wire n_797, n_800, n_802, n_803, n_806, n_808, n_811, n_814;
  wire n_819, n_821, n_823, n_828, n_832, n_834, n_846, n_848;
  wire n_850, n_852, n_853, n_854, n_855, n_857, n_858, n_859;
  wire n_860, n_861, n_863, n_864, n_865, n_866, n_869, n_871;
  wire n_872, n_875, n_878, n_880, n_883, n_889, n_894, n_898;
  wire n_900, n_914, n_915, n_918, n_920, n_921, n_922, n_923;
  wire n_925, n_926, n_927, n_928, n_929, n_931, n_932, n_933;
  wire n_935, n_937, n_938, n_941, n_943, n_944, n_947, n_949;
  wire n_954, n_957, n_962, n_966, n_971, n_975, n_977, n_998;
  wire n_1000, n_1001, n_1002, n_1003, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1011, n_1012, n_1013, n_1015, n_1017, n_1018, n_1021;
  wire n_1023, n_1024, n_1027, n_1029, n_1034, n_1037, n_1042, n_1047;
  wire n_1054, n_1058, n_1060, n_1075, n_1077, n_1079, n_1081, n_1082;
  wire n_1083, n_1084, n_1086, n_1087, n_1088, n_1089, n_1090, n_1092;
  wire n_1093, n_1094, n_1095, n_1098, n_1100, n_1101, n_1104, n_1107;
  wire n_1109, n_1112, n_1118, n_1123, n_1127, n_1129, n_1143, n_1144;
  wire n_1147, n_1149, n_1150, n_1151, n_1152, n_1154, n_1155, n_1156;
  wire n_1157, n_1158, n_1160, n_1161, n_1162, n_1164, n_1166, n_1167;
  wire n_1170, n_1172, n_1173, n_1176, n_1178, n_1183, n_1186, n_1191;
  wire n_1195, n_1200, n_1204, n_1206, n_1227, n_1229, n_1230, n_1231;
  wire n_1232, n_1234, n_1235, n_1236, n_1237, n_1238, n_1240, n_1241;
  wire n_1242, n_1244, n_1246, n_1247, n_1250, n_1252, n_1253, n_1256;
  wire n_1258, n_1263, n_1266, n_1271, n_1276, n_1283, n_1287, n_1289;
  wire n_1304, n_1306, n_1308, n_1310, n_1311, n_1312, n_1313, n_1315;
  wire n_1316, n_1317, n_1318, n_1319, n_1321, n_1322, n_1323, n_1324;
  wire n_1327, n_1329, n_1330, n_1333, n_1336, n_1338, n_1341, n_1347;
  wire n_1352, n_1356, n_1358, n_1372, n_1373, n_1376, n_1378, n_1379;
  wire n_1380, n_1381, n_1383, n_1384, n_1385, n_1386, n_1387, n_1389;
  wire n_1390, n_1391, n_1393, n_1395, n_1396, n_1399, n_1401, n_1402;
  wire n_1405, n_1407, n_1412, n_1415, n_1420, n_1424, n_1429, n_1433;
  wire n_1435, n_1456, n_1458, n_1459, n_1460, n_1461, n_1463, n_1464;
  wire n_1465, n_1466, n_1467, n_1469, n_1470, n_1471, n_1473, n_1475;
  wire n_1476, n_1479, n_1481, n_1482, n_1485, n_1487, n_1492, n_1495;
  wire n_1500, n_1505, n_1512, n_1516, n_1518, n_1535, n_1540, n_1542;
  wire n_1546, n_1548, n_1552, n_1553, n_1556, n_1558, n_1562, n_1565;
  wire n_1567, n_1576, n_1608, n_1610, n_1614, n_1616, n_1620, n_1622;
  wire n_1625, n_1628, n_1630, n_1634, n_1636, n_1641, n_1649, n_1653;
  wire n_1688, n_1690, n_1694, n_1696, n_1700, n_1702, n_1705, n_1708;
  wire n_1710, n_1714, n_1716, n_1721, n_1729, n_1734, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815;
  wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  wire n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1840;
  wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1865, n_1866;
  wire n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874;
  wire n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882;
  wire n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890;
  wire n_1891, n_1892, n_1893, n_1894, n_1895, n_1898, n_1899, n_1900;
  wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908;
  wire n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916;
  wire n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924;
  wire n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932;
  wire n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1940, n_1941;
  wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
  wire n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957;
  wire n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965;
  wire n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973;
  wire n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1982;
  wire n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990;
  wire n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998;
  wire n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006;
  wire n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014;
  wire n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022;
  wire n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031;
  wire n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039;
  wire n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047;
  wire n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
  wire n_2072;
  not g1 (QUOTIENT[14], n_39);
  nand g11 (QUOTIENT[13], n_56, n_59);
  and g19 (n_82, n_535, n_81);
  and g31 (n_112, n_709, n_111);
  or g46 (QUOTIENT[6], n_151, n_147);
  or g58 (QUOTIENT[4], n_196, n_192);
  or g70 (QUOTIENT[2], n_241, n_237);
  or g82 (QUOTIENT[0], n_286, n_2072);
  xor g84 (n_349, B[0], B[1]);
  nand g2 (n_302, B[0], B[1]);
  nor g87 (n_305, B[1], B[2]);
  nand g88 (n_308, B[1], B[2]);
  nand g90 (n_310, B[2], B[3]);
  nand g92 (n_312, B[3], B[4]);
  nand g13 (n_316, B[4], B[5]);
  nand g15 (n_318, B[5], B[6]);
  nand g95 (n_322, n_308, n_1779);
  nor g96 (n_313, n_310, n_311);
  nor g24 (n_325, n_358, n_311);
  nor g25 (n_319, n_316, n_317);
  nor g99 (n_331, n_360, n_317);
  nand g102 (n_342, n_310, n_1816);
  nand g103 (n_327, n_325, n_322);
  nand g104 (n_332, n_1783, n_327);
  nand g38 (n_336, n_331, B[6]);
  nand g107 (n_346, n_316, n_1829);
  nand g108 (n_335, n_331, n_332);
  nand g109 (n_348, n_329, n_335);
  xnor g50 (n_42, n_322, n_1780);
  xnor g115 (n_43, n_342, n_1782);
  xnor g117 (n_44, n_332, n_1784);
  xnor g120 (n_45, n_346, n_1785);
  nor g126 (n_358, B[2], B[3]);
  nor g36 (n_360, B[4], B[5]);
  nand g158 (n_384, n_379, n_1793);
  nor g159 (n_382, n_381, B[3]);
  nor g160 (n_387, n_383, B[3]);
  nand g165 (n_388, n_387, n_384);
  xnor g175 (n_49, n_377, n_1796);
  xnor g177 (n_51, n_384, n_1832);
  nand g197 (n_416, n_411, n_408);
  nor g198 (n_414, n_413, B[2]);
  nor g199 (n_419, n_415, B[2]);
  nor g200 (n_311, B[3], B[4]);
  nor g201 (n_317, B[5], B[6]);
  nand g205 (n_420, n_419, n_416);
  nand g209 (n_431, n_311, n_317);
  xnor g220 (n_52, n_416, n_1833);
  nand g243 (n_453, n_448, n_1815);
  nor g244 (n_451, n_450, n_42);
  nor g245 (n_456, n_452, n_42);
  nor g246 (n_458, n_43, n_44);
  nor g247 (n_460, n_45, n_46);
  nand g251 (n_457, n_456, n_453);
  nand g255 (n_468, n_458, n_460);
  xnor g266 (n_50, n_377, n_1817);
  xnor g268 (n_53, n_453, n_1834);
  nand g303 (n_502, n_491, n_1798);
  nor g304 (n_496, n_493, n_494);
  nor g307 (n_505, n_498, n_494);
  nor g308 (n_500, n_499, B[5]);
  nor g309 (n_510, n_501, B[5]);
  nand g312 (n_522, n_493, n_1850);
  nand g313 (n_507, n_505, n_502);
  nand g314 (n_512, n_1840, n_507);
  xnor g327 (n_67, n_489, n_1799);
  xnor g329 (n_69, n_502, n_1847);
  xnor g332 (n_72, n_522, n_1851);
  xnor g334 (n_75, n_512, n_1844);
  nand g359 (n_550, n_539, n_536);
  nor g360 (n_544, n_541, n_542);
  nor g363 (n_553, n_546, n_542);
  nor g364 (n_548, n_547, B[4]);
  nor g365 (n_558, n_549, B[4]);
  nand g369 (n_576, n_541, n_1852);
  nand g370 (n_555, n_553, n_550);
  nand g371 (n_563, n_1842, n_555);
  nand g377 (n_570, n_558, n_317);
  xnor g392 (n_70, n_550, n_1848);
  xnor g395 (n_73, n_576, n_1853);
  xnor g397 (n_76, n_563, n_1845);
  nand g423 (n_605, n_594, n_1818);
  nor g424 (n_599, n_596, n_597);
  nor g427 (n_608, n_601, n_597);
  nor g428 (n_603, n_602, n_44);
  nor g429 (n_613, n_604, n_44);
  nand g433 (n_633, n_596, n_1854);
  nand g434 (n_610, n_608, n_605);
  nand g435 (n_618, n_1843, n_610);
  nand g441 (n_625, n_613, n_460);
  xnor g456 (n_68, n_489, n_1819);
  xnor g458 (n_71, n_605, n_1849);
  xnor g461 (n_74, n_633, n_1855);
  xnor g463 (n_77, n_618, n_1846);
  nand g502 (n_668, n_654, n_1801);
  nor g503 (n_659, n_656, n_657);
  nor g506 (n_671, n_661, n_657);
  nor g507 (n_665, n_662, n_663);
  nor g510 (n_679, n_667, n_663);
  nand g513 (n_692, n_656, n_1875);
  nand g514 (n_673, n_671, n_668);
  nand g515 (n_681, n_1865, n_673);
  nor g516 (n_677, n_674, n_675);
  nand g523 (n_696, n_662, n_1893);
  nand g524 (n_684, n_679, n_681);
  nand g525 (n_698, n_675, n_684);
  nand g528 (n_650, n_1889, n_1890);
  xnor g530 (n_91, n_652, n_1802);
  xnor g532 (n_93, n_668, n_1872);
  xnor g535 (n_96, n_692, n_1876);
  xnor g537 (n_99, n_681, n_1881);
  xnor g540 (n_102, n_696, n_1884);
  xnor g542 (n_105, n_698, n_1869);
  nand g569 (n_730, n_713, n_710);
  nor g570 (n_718, n_715, n_716);
  nor g573 (n_733, n_720, n_716);
  nor g574 (n_724, n_721, n_722);
  nor g577 (n_739, n_726, n_722);
  nor g578 (n_728, n_727, B[6]);
  nor g579 (n_741, n_729, B[6]);
  nand g582 (n_759, n_715, n_1877);
  nand g583 (n_735, n_733, n_730);
  nand g584 (n_744, n_1867, n_735);
  nor g592 (n_754, n_1887, n_728);
  nand g593 (n_752, n_739, n_741);
  nand g596 (n_763, n_721, n_1894);
  nand g597 (n_747, n_739, n_744);
  nand g598 (n_765, n_736, n_747);
  nand g604 (n_709, n_754, n_1891);
  xnor g608 (n_94, n_730, n_1873);
  xnor g611 (n_97, n_759, n_1878);
  xnor g613 (n_100, n_744, n_1882);
  xnor g616 (n_103, n_763, n_1885);
  xnor g618 (n_106, n_765, n_1870);
  nand g645 (n_797, n_780, n_1820);
  nor g646 (n_785, n_782, n_783);
  nor g649 (n_800, n_787, n_783);
  nor g650 (n_791, n_788, n_789);
  nor g653 (n_806, n_793, n_789);
  nor g654 (n_795, n_794, n_46);
  nor g655 (n_808, n_796, n_46);
  nand g658 (n_828, n_782, n_1879);
  nand g659 (n_802, n_800, n_797);
  nand g660 (n_811, n_1868, n_802);
  nor g668 (n_821, n_1888, n_795);
  nand g669 (n_819, n_806, n_808);
  nand g672 (n_832, n_788, n_1895);
  nand g673 (n_814, n_806, n_811);
  nand g674 (n_834, n_803, n_814);
  nand g680 (n_823, n_821, n_1892);
  xnor g684 (n_92, n_652, n_1821);
  xnor g686 (n_95, n_797, n_1874);
  xnor g689 (n_98, n_828, n_1880);
  xnor g691 (n_101, n_811, n_1883);
  xnor g694 (n_104, n_832, n_1886);
  xnor g696 (n_107, n_834, n_1871);
  nand g732 (n_866, n_850, n_1804);
  nor g733 (n_855, n_852, n_853);
  nor g736 (n_869, n_857, n_853);
  nor g737 (n_861, n_858, n_859);
  nor g740 (n_875, n_863, n_859);
  nand g744 (n_894, n_852, n_1915);
  nand g745 (n_871, n_869, n_866);
  nand g746 (n_880, n_1903, n_871);
  nor g751 (n_878, n_872, n_865);
  nand g757 (n_898, n_858, n_1935);
  nand g758 (n_883, n_875, n_880);
  nand g759 (n_900, n_872, n_883);
  nand g763 (n_889, n_1929, n_1930);
  xnor g766 (n_123, n_848, n_1805);
  xnor g768 (n_125, n_866, n_1912);
  xnor g771 (n_128, n_894, n_1916);
  xnor g773 (n_131, n_880, n_1921);
  xnor g776 (n_134, n_898, n_1924);
  xnor g778 (n_137, n_900, n_1909);
  nand g812 (n_938, n_918, n_915);
  nor g813 (n_923, n_920, n_921);
  nor g816 (n_941, n_925, n_921);
  nor g817 (n_929, n_926, n_927);
  nor g820 (n_947, n_931, n_927);
  nor g821 (n_935, n_932, n_933);
  nor g824 (n_949, n_937, n_933);
  nand g827 (n_971, n_920, n_1917);
  nand g828 (n_943, n_941, n_938);
  nand g829 (n_954, n_1906, n_943);
  nand g839 (n_962, n_947, n_949);
  nand g842 (n_975, n_926, n_1936);
  nand g843 (n_957, n_947, n_954);
  nand g844 (n_977, n_944, n_957);
  nand g850 (n_966, n_1931, n_1932);
  xnor g855 (n_126, n_938, n_1913);
  xnor g858 (n_129, n_971, n_1918);
  xnor g860 (n_132, n_954, n_1922);
  xnor g863 (n_135, n_975, n_1925);
  xnor g865 (n_138, n_977, n_1910);
  nand g904 (n_1018, n_998, n_1822);
  nor g905 (n_1003, n_1000, n_1001);
  nor g908 (n_1021, n_1005, n_1001);
  nor g909 (n_1009, n_1006, n_1007);
  nor g912 (n_1027, n_1011, n_1007);
  nor g913 (n_1015, n_1012, n_1013);
  nor g916 (n_1029, n_1017, n_1013);
  nand g919 (n_1054, n_1000, n_1919);
  nand g920 (n_1023, n_1021, n_1018);
  nand g921 (n_1034, n_1908, n_1023);
  nand g931 (n_1042, n_1027, n_1029);
  nand g934 (n_1058, n_1006, n_1937);
  nand g935 (n_1037, n_1027, n_1034);
  nand g936 (n_1060, n_1024, n_1037);
  nand g942 (n_1047, n_1933, n_1934);
  nand g945 (n_151, n_1899, n_1938);
  xnor g947 (n_124, n_848, n_1823);
  xnor g949 (n_127, n_1018, n_1914);
  xnor g952 (n_130, n_1054, n_1920);
  xnor g954 (n_133, n_1034, n_1923);
  xnor g957 (n_136, n_1058, n_1926);
  xnor g959 (n_139, n_1060, n_1911);
  nand g1000 (n_1095, n_1079, n_1807);
  nor g1001 (n_1084, n_1081, n_1082);
  nor g1004 (n_1098, n_1086, n_1082);
  nor g1005 (n_1090, n_1087, n_1088);
  nor g1008 (n_1104, n_1092, n_1088);
  nand g1012 (n_1123, n_1081, n_1957);
  nand g1013 (n_1100, n_1098, n_1095);
  nand g1014 (n_1109, n_1945, n_1100);
  nor g1019 (n_1107, n_1101, n_1094);
  nand g1025 (n_1127, n_1087, n_1977);
  nand g1026 (n_1112, n_1104, n_1109);
  nand g1027 (n_1129, n_1101, n_1112);
  nand g1031 (n_1118, n_1971, n_1972);
  xnor g1034 (n_165, n_1077, n_1808);
  xnor g1036 (n_168, n_1095, n_1954);
  xnor g1039 (n_171, n_1123, n_1958);
  xnor g1041 (n_174, n_1109, n_1963);
  xnor g1044 (n_177, n_1127, n_1966);
  xnor g1046 (n_180, n_1129, n_1951);
  nand g1080 (n_1167, n_1147, n_1144);
  nor g1081 (n_1152, n_1149, n_1150);
  nor g1084 (n_1170, n_1154, n_1150);
  nor g1085 (n_1158, n_1155, n_1156);
  nor g1088 (n_1176, n_1160, n_1156);
  nor g1089 (n_1164, n_1161, n_1162);
  nor g1092 (n_1178, n_1166, n_1162);
  nand g1095 (n_1200, n_1149, n_1959);
  nand g1096 (n_1172, n_1170, n_1167);
  nand g1097 (n_1183, n_1948, n_1172);
  nand g1107 (n_1191, n_1176, n_1178);
  nand g1110 (n_1204, n_1155, n_1978);
  nand g1111 (n_1186, n_1176, n_1183);
  nand g1112 (n_1206, n_1173, n_1186);
  nand g1118 (n_1195, n_1973, n_1974);
  xnor g1123 (n_169, n_1167, n_1955);
  xnor g1126 (n_172, n_1200, n_1960);
  xnor g1128 (n_175, n_1183, n_1964);
  xnor g1131 (n_178, n_1204, n_1967);
  xnor g1133 (n_181, n_1206, n_1952);
  nand g1172 (n_1247, n_1227, n_1824);
  nor g1173 (n_1232, n_1229, n_1230);
  nor g1176 (n_1250, n_1234, n_1230);
  nor g1177 (n_1238, n_1235, n_1236);
  nor g1180 (n_1256, n_1240, n_1236);
  nor g1181 (n_1244, n_1241, n_1242);
  nor g1184 (n_1258, n_1246, n_1242);
  nand g1187 (n_1283, n_1229, n_1961);
  nand g1188 (n_1252, n_1250, n_1247);
  nand g1189 (n_1263, n_1950, n_1252);
  nand g1199 (n_1271, n_1256, n_1258);
  nand g1202 (n_1287, n_1235, n_1979);
  nand g1203 (n_1266, n_1256, n_1263);
  nand g1204 (n_1289, n_1253, n_1266);
  nand g1210 (n_1276, n_1975, n_1976);
  nand g1213 (n_196, n_1941, n_1980);
  xnor g1215 (n_167, n_1077, n_1825);
  xnor g1217 (n_170, n_1247, n_1956);
  xnor g1220 (n_173, n_1283, n_1962);
  xnor g1222 (n_176, n_1263, n_1965);
  xnor g1225 (n_179, n_1287, n_1968);
  xnor g1227 (n_182, n_1289, n_1953);
  nand g1268 (n_1324, n_1308, n_1810);
  nor g1269 (n_1313, n_1310, n_1311);
  nor g1272 (n_1327, n_1315, n_1311);
  nor g1273 (n_1319, n_1316, n_1317);
  nor g1276 (n_1333, n_1321, n_1317);
  nand g1280 (n_1352, n_1310, n_1999);
  nand g1281 (n_1329, n_1327, n_1324);
  nand g1282 (n_1338, n_1987, n_1329);
  nor g1287 (n_1336, n_1330, n_1323);
  nand g1293 (n_1356, n_1316, n_2019);
  nand g1294 (n_1341, n_1333, n_1338);
  nand g1295 (n_1358, n_1330, n_1341);
  nand g1299 (n_1347, n_2013, n_2014);
  xnor g1302 (n_210, n_1306, n_1811);
  xnor g1304 (n_213, n_1324, n_1996);
  xnor g1307 (n_216, n_1352, n_2000);
  xnor g1309 (n_219, n_1338, n_2005);
  xnor g1312 (n_222, n_1356, n_2008);
  xnor g1314 (n_225, n_1358, n_1993);
  nand g1348 (n_1396, n_1376, n_1373);
  nor g1349 (n_1381, n_1378, n_1379);
  nor g1352 (n_1399, n_1383, n_1379);
  nor g1353 (n_1387, n_1384, n_1385);
  nor g1356 (n_1405, n_1389, n_1385);
  nor g1357 (n_1393, n_1390, n_1391);
  nor g1360 (n_1407, n_1395, n_1391);
  nand g1363 (n_1429, n_1378, n_2001);
  nand g1364 (n_1401, n_1399, n_1396);
  nand g1365 (n_1412, n_1990, n_1401);
  nand g1375 (n_1420, n_1405, n_1407);
  nand g1378 (n_1433, n_1384, n_2020);
  nand g1379 (n_1415, n_1405, n_1412);
  nand g1380 (n_1435, n_1402, n_1415);
  nand g1386 (n_1424, n_2015, n_2016);
  xnor g1391 (n_214, n_1396, n_1997);
  xnor g1394 (n_217, n_1429, n_2002);
  xnor g1396 (n_220, n_1412, n_2006);
  xnor g1399 (n_223, n_1433, n_2009);
  xnor g1401 (n_226, n_1435, n_1994);
  nand g1440 (n_1476, n_1456, n_1826);
  nor g1441 (n_1461, n_1458, n_1459);
  nor g1444 (n_1479, n_1463, n_1459);
  nor g1445 (n_1467, n_1464, n_1465);
  nor g1448 (n_1485, n_1469, n_1465);
  nor g1449 (n_1473, n_1470, n_1471);
  nor g1452 (n_1487, n_1475, n_1471);
  nand g1455 (n_1512, n_1458, n_2003);
  nand g1456 (n_1481, n_1479, n_1476);
  nand g1457 (n_1492, n_1992, n_1481);
  nand g1467 (n_1500, n_1485, n_1487);
  nand g1470 (n_1516, n_1464, n_2021);
  nand g1471 (n_1495, n_1485, n_1492);
  nand g1472 (n_1518, n_1482, n_1495);
  nand g1478 (n_1505, n_2017, n_2018);
  nand g1481 (n_241, n_1983, n_2022);
  xnor g1483 (n_212, n_1306, n_1827);
  xnor g1485 (n_215, n_1476, n_1998);
  xnor g1488 (n_218, n_1512, n_2004);
  xnor g1490 (n_221, n_1492, n_2007);
  xnor g1493 (n_224, n_1516, n_2010);
  xnor g1495 (n_227, n_1518, n_1995);
  nand g1536 (n_1553, n_1775, n_1813);
  nor g1537 (n_1542, n_2036, n_1540);
  nor g1540 (n_1556, n_2038, n_1540);
  nor g1541 (n_1548, n_2033, n_1546);
  nor g1544 (n_1562, n_2039, n_1546);
  nand g1549 (n_1558, n_1556, n_1553);
  nand g1550 (n_1567, n_2056, n_1558);
  nor g1555 (n_1565, n_2054, n_1552);
  nand g1567 (n_1576, n_2065, n_2066);
  nand g1616 (n_1625, n_1773, n_1774);
  nor g1617 (n_1610, n_2029, n_1608);
  nor g1620 (n_1628, n_2031, n_1608);
  nor g1621 (n_1616, n_2024, n_1614);
  nor g1624 (n_1634, n_2032, n_1614);
  nor g1625 (n_1622, n_2027, n_1620);
  nor g1628 (n_1636, n_2026, n_1620);
  nand g1632 (n_1630, n_1628, n_1625);
  nand g1633 (n_1641, n_2053, n_1630);
  nand g1643 (n_1649, n_1634, n_1636);
  nand g1654 (n_1653, n_2063, n_2064);
  nand g1708 (n_1705, n_1791, n_1828);
  nor g1709 (n_1690, n_2046, n_1688);
  nor g1712 (n_1708, n_2048, n_1688);
  nor g1713 (n_1696, n_2041, n_1694);
  nor g1716 (n_1714, n_2049, n_1694);
  nor g1717 (n_1702, n_2044, n_1700);
  nor g1720 (n_1716, n_2043, n_1700);
  nand g1724 (n_1710, n_1708, n_1705);
  nand g1725 (n_1721, n_2060, n_1710);
  nand g1735 (n_1729, n_1714, n_1716);
  nand g1746 (n_1734, n_2067, n_2068);
  nand g1749 (n_286, n_2040, n_2069);
  or g1781 (n_1758, wc, A[14]);
  not gc (wc, B[0]);
  or g1782 (n_1759, B[6], wc0);
  not gc0 (wc0, n_360);
  xnor g1783 (n_1760, A[14], B[0]);
  or g1784 (n_379, B[1], wc1);
  not gc1 (wc1, A[13]);
  or g1785 (n_377, wc2, A[12]);
  not gc2 (wc2, B[0]);
  and g1786 (n_1761, B[1], wc3);
  not gc3 (wc3, A[13]);
  or g1787 (n_411, B[0], wc4);
  not gc4 (wc4, A[13]);
  and g1788 (n_408, B[0], wc5);
  not gc5 (wc5, A[13]);
  xnor g1789 (n_1762, A[12], B[0]);
  or g1790 (n_491, B[1], wc6);
  not gc6 (wc6, A[11]);
  or g1791 (n_489, wc7, A[10]);
  not gc7 (wc7, B[0]);
  and g1792 (n_1763, B[1], wc8);
  not gc8 (wc8, A[11]);
  or g1793 (n_539, B[0], wc9);
  not gc9 (wc9, A[11]);
  and g1794 (n_536, B[0], wc10);
  not gc10 (wc10, A[11]);
  xnor g1795 (n_1764, A[10], B[0]);
  or g1796 (n_654, B[1], wc11);
  not gc11 (wc11, A[9]);
  or g1797 (n_652, wc12, A[8]);
  not gc12 (wc12, B[0]);
  and g1798 (n_1765, B[1], wc13);
  not gc13 (wc13, A[9]);
  or g1799 (n_713, B[0], wc14);
  not gc14 (wc14, A[9]);
  and g1800 (n_710, B[0], wc15);
  not gc15 (wc15, A[9]);
  xnor g1801 (n_1766, A[8], B[0]);
  or g1802 (n_850, B[1], wc16);
  not gc16 (wc16, A[7]);
  or g1803 (n_848, wc17, A[6]);
  not gc17 (wc17, B[0]);
  and g1804 (n_1767, B[1], wc18);
  not gc18 (wc18, A[7]);
  or g1805 (n_918, B[0], wc19);
  not gc19 (wc19, A[7]);
  and g1806 (n_915, B[0], wc20);
  not gc20 (wc20, A[7]);
  xnor g1807 (n_1768, A[6], B[0]);
  or g1808 (n_1079, B[1], wc21);
  not gc21 (wc21, A[5]);
  or g1809 (n_1077, wc22, A[4]);
  not gc22 (wc22, B[0]);
  and g1810 (n_1769, B[1], wc23);
  not gc23 (wc23, A[5]);
  or g1811 (n_1147, B[0], wc24);
  not gc24 (wc24, A[5]);
  and g1812 (n_1144, B[0], wc25);
  not gc25 (wc25, A[5]);
  xnor g1813 (n_1770, A[4], B[0]);
  or g1814 (n_1308, B[1], wc26);
  not gc26 (wc26, A[3]);
  or g1815 (n_1306, wc27, A[2]);
  not gc27 (wc27, B[0]);
  and g1816 (n_1771, B[1], wc28);
  not gc28 (wc28, A[3]);
  or g1817 (n_1376, B[0], wc29);
  not gc29 (wc29, A[3]);
  and g1818 (n_1373, B[0], wc30);
  not gc30 (wc30, A[3]);
  xnor g1819 (n_1772, A[2], B[0]);
  or g1820 (n_1773, B[0], wc31);
  not gc31 (wc31, A[1]);
  and g1821 (n_1774, B[0], wc32);
  not gc32 (wc32, A[1]);
  or g1822 (n_1775, B[1], wc33);
  not gc33 (wc33, A[1]);
  or g1823 (n_1535, wc34, A[0]);
  not gc34 (wc34, B[0]);
  and g1824 (n_1776, B[1], wc35);
  not gc35 (wc35, A[1]);
  or g1825 (n_1777, B[1], wc36);
  not gc36 (wc36, n_1758);
  or g1826 (n_1778, wc37, n_305);
  not gc37 (wc37, n_308);
  or g1827 (n_1779, n_302, n_305);
  or g1828 (n_1780, n_358, wc38);
  not gc38 (wc38, n_310);
  or g1829 (n_448, wc39, n_349);
  not gc39 (wc39, A[13]);
  and g1830 (n_1781, wc40, n_349);
  not gc40 (wc40, A[13]);
  or g1831 (n_1782, n_311, wc41);
  not gc41 (wc41, n_312);
  and g1832 (n_1783, wc42, n_312);
  not gc42 (wc42, n_313);
  or g1833 (n_1784, n_360, wc43);
  not gc43 (wc43, n_316);
  or g1834 (n_1785, n_317, wc44);
  not gc44 (wc44, n_318);
  and g1835 (n_329, wc45, n_318);
  not gc45 (wc45, n_319);
  or g1836 (n_594, wc46, n_349);
  not gc46 (wc46, A[11]);
  and g1837 (n_1786, wc47, n_349);
  not gc47 (wc47, A[11]);
  or g1838 (n_780, wc48, n_349);
  not gc48 (wc48, A[9]);
  and g1839 (n_1787, wc49, n_349);
  not gc49 (wc49, A[9]);
  or g1840 (n_998, wc50, n_349);
  not gc50 (wc50, A[7]);
  and g1841 (n_1788, wc51, n_349);
  not gc51 (wc51, A[7]);
  or g1842 (n_1227, wc52, n_349);
  not gc52 (wc52, A[5]);
  and g1843 (n_1789, wc53, n_349);
  not gc53 (wc53, A[5]);
  or g1844 (n_1456, wc54, n_349);
  not gc54 (wc54, A[3]);
  and g1845 (n_1790, wc55, n_349);
  not gc55 (wc55, A[3]);
  or g1846 (n_1791, wc56, n_349);
  not gc56 (wc56, A[1]);
  and g1847 (n_1792, wc57, n_349);
  not gc57 (wc57, A[1]);
  or g1848 (n_1793, n_1761, wc58);
  not gc58 (wc58, n_377);
  xor g1849 (n_1794, n_302, n_1778);
  and g1850 (n_1795, B[6], wc59);
  not gc59 (wc59, n_329);
  or g1851 (n_1796, n_1761, wc60);
  not gc60 (wc60, n_379);
  or g1852 (n_1797, n_408, wc61);
  not gc61 (wc61, n_411);
  or g1853 (n_1798, n_1763, wc62);
  not gc62 (wc62, n_489);
  or g1854 (n_1799, n_1763, wc63);
  not gc63 (wc63, n_491);
  or g1855 (n_1800, n_536, wc64);
  not gc64 (wc64, n_539);
  or g1856 (n_1801, n_1765, wc65);
  not gc65 (wc65, n_652);
  or g1857 (n_1802, n_1765, wc66);
  not gc66 (wc66, n_654);
  or g1858 (n_1803, n_710, wc67);
  not gc67 (wc67, n_713);
  or g1859 (n_1804, n_1767, wc68);
  not gc68 (wc68, n_848);
  or g1860 (n_1805, n_1767, wc69);
  not gc69 (wc69, n_850);
  or g1861 (n_1806, n_915, wc70);
  not gc70 (wc70, n_918);
  or g1862 (n_1807, n_1769, wc71);
  not gc71 (wc71, n_1077);
  or g1863 (n_1808, n_1769, wc72);
  not gc72 (wc72, n_1079);
  or g1864 (n_1809, n_1144, wc73);
  not gc73 (wc73, n_1147);
  or g1865 (n_1810, n_1771, wc74);
  not gc74 (wc74, n_1306);
  or g1866 (n_1811, n_1771, wc75);
  not gc75 (wc75, n_1308);
  or g1867 (n_1812, n_1373, wc76);
  not gc76 (wc76, n_1376);
  or g1868 (n_1813, n_1776, wc77);
  not gc77 (wc77, n_1535);
  or g1869 (n_1814, n_1777, wc78);
  not gc78 (wc78, n_358);
  or g1870 (n_1815, n_1781, wc79);
  not gc79 (wc79, n_377);
  or g1871 (n_1816, n_358, wc80);
  not gc80 (wc80, n_322);
  or g1872 (n_1817, n_1781, wc81);
  not gc81 (wc81, n_448);
  or g1873 (n_1818, n_1786, wc82);
  not gc82 (wc82, n_489);
  or g1874 (n_1819, n_1786, wc83);
  not gc83 (wc83, n_594);
  or g1875 (n_1820, n_1787, wc84);
  not gc84 (wc84, n_652);
  or g1876 (n_1821, n_1787, wc85);
  not gc85 (wc85, n_780);
  or g1877 (n_1822, n_1788, wc86);
  not gc86 (wc86, n_848);
  or g1878 (n_1823, n_1788, wc87);
  not gc87 (wc87, n_998);
  or g1879 (n_1824, n_1789, wc88);
  not gc88 (wc88, n_1077);
  or g1880 (n_1825, n_1789, wc89);
  not gc89 (wc89, n_1227);
  or g1881 (n_1826, n_1790, wc90);
  not gc90 (wc90, n_1306);
  or g1882 (n_1827, n_1790, wc91);
  not gc91 (wc91, n_1456);
  or g1883 (n_1828, n_1792, wc92);
  not gc92 (wc92, n_1535);
  or g1884 (n_39, n_1759, n_1814);
  or g1885 (n_1829, n_360, wc93);
  not gc93 (wc93, n_332);
  or g1886 (n_1830, n_336, wc94);
  not gc94 (wc94, n_332);
  or g1887 (n_1831, wc95, n_1795);
  not gc95 (wc95, n_1830);
  or g1888 (n_40, wc96, wc99);
  and gc99 (wc99, A[14], n_39);
  and gc98 (wc96, wc97, wc98);
  not gc97 (wc98, n_1760);
  not gc96 (wc97, n_39);
  xor g1889 (n_46, n_348, B[6]);
  or g1890 (n_381, B[2], wc100);
  not gc100 (wc100, n_40);
  and g1891 (n_383, B[2], wc101);
  not gc101 (wc101, n_40);
  or g1892 (n_413, B[1], wc102);
  not gc102 (wc102, n_40);
  and g1893 (n_415, B[1], wc103);
  not gc103 (wc103, n_40);
  or g1894 (n_450, wc104, n_1794);
  not gc104 (wc104, n_40);
  and g1895 (n_452, wc105, n_1794);
  not gc105 (wc105, n_40);
  or g1896 (n_1832, n_383, wc106);
  not gc106 (wc106, n_381);
  or g1897 (n_1833, n_415, wc107);
  not gc107 (wc107, n_413);
  or g1898 (n_1834, n_452, wc108);
  not gc108 (wc108, n_450);
  or g1899 (n_1835, wc109, n_382);
  not gc109 (wc109, n_388);
  or g1900 (n_1836, wc110, n_414);
  not gc110 (wc110, n_420);
  or g1901 (n_1837, wc111, n_451);
  not gc111 (wc111, n_457);
  or g1902 (n_54, wc112, n_1759);
  not gc112 (wc112, n_1835);
  or g1903 (n_56, wc113, n_431);
  not gc113 (wc113, n_1836);
  or g1904 (n_1838, wc114, n_468);
  not gc114 (wc114, n_1837);
  and g1905 (n_57, n_56, wc115);
  not gc115 (wc115, n_54);
  or g1906 (n_59, n_1831, n_1838);
  and g1907 (n_60, n_59, wc116);
  not gc116 (wc116, n_56);
  or g1908 (QUOTIENT[12], wc117, n_57);
  not gc117 (wc117, n_59);
  or g1909 (n_65, wc118, wc119, wc120, wc121);
  and gc122 (wc121, wc122, n_53);
  not gc121 (wc122, n_59);
  and gc120 (wc120, n_60, n_52);
  and gc119 (wc119, n_57, n_51);
  and gc118 (wc118, n_54, n_40);
  or g1910 (n_63, wc123, wc124, wc126, wc127);
  and gc129 (wc127, wc128, wc129);
  not gc128 (wc129, n_1762);
  not gc127 (wc128, n_59);
  and gc126 (wc126, A[12], n_60);
  and gc125 (wc124, n_57, wc125);
  not gc124 (wc125, n_1762);
  and gc123 (wc123, A[12], n_54);
  or g1911 (n_64, wc130, wc131, wc132, wc133);
  and gc134 (wc133, wc134, n_50);
  not gc133 (wc134, n_59);
  and gc132 (wc132, n_60, n_1797);
  and gc131 (wc131, n_57, n_49);
  and gc130 (wc130, A[13], n_54);
  or g1912 (n_499, B[4], wc135);
  not gc135 (wc135, n_65);
  or g1913 (n_493, B[2], wc136);
  not gc136 (wc136, n_63);
  and g1914 (n_494, B[3], wc137);
  not gc137 (wc137, n_64);
  or g1915 (n_495, B[3], wc138);
  not gc138 (wc138, n_64);
  and g1916 (n_498, B[2], wc139);
  not gc139 (wc139, n_63);
  and g1917 (n_501, B[4], wc140);
  not gc140 (wc140, n_65);
  or g1918 (n_547, B[3], wc141);
  not gc141 (wc141, n_65);
  or g1919 (n_541, B[1], wc142);
  not gc142 (wc142, n_63);
  and g1920 (n_542, B[2], wc143);
  not gc143 (wc143, n_64);
  or g1921 (n_543, B[2], wc144);
  not gc144 (wc144, n_64);
  and g1922 (n_546, B[1], wc145);
  not gc145 (wc145, n_63);
  and g1923 (n_549, B[3], wc146);
  not gc146 (wc146, n_65);
  or g1924 (n_602, wc147, n_43);
  not gc147 (wc147, n_65);
  or g1925 (n_596, wc148, n_1794);
  not gc148 (wc148, n_63);
  and g1926 (n_597, wc149, n_42);
  not gc149 (wc149, n_64);
  or g1927 (n_598, wc150, n_42);
  not gc150 (wc150, n_64);
  and g1928 (n_601, wc151, n_1794);
  not gc151 (wc151, n_63);
  and g1929 (n_604, wc152, n_43);
  not gc152 (wc152, n_65);
  and g1930 (n_1840, n_495, wc153);
  not gc153 (wc153, n_496);
  or g1931 (n_1841, B[6], wc154);
  not gc154 (wc154, n_510);
  and g1932 (n_1842, n_543, wc155);
  not gc155 (wc155, n_544);
  and g1933 (n_1843, n_598, wc156);
  not gc156 (wc156, n_599);
  or g1934 (n_1844, n_501, wc157);
  not gc157 (wc157, n_499);
  or g1935 (n_1845, n_549, wc158);
  not gc158 (wc158, n_547);
  or g1936 (n_1846, n_604, wc159);
  not gc159 (wc159, n_602);
  or g1937 (n_1847, n_498, wc160);
  not gc160 (wc160, n_493);
  or g1938 (n_1848, n_546, wc161);
  not gc161 (wc161, n_541);
  or g1939 (n_1849, n_601, wc162);
  not gc162 (wc162, n_596);
  or g1940 (n_1850, n_498, wc163);
  not gc163 (wc163, n_502);
  or g1941 (n_1851, wc164, n_494);
  not gc164 (wc164, n_495);
  or g1942 (n_1852, n_546, wc165);
  not gc165 (wc165, n_550);
  or g1943 (n_1853, wc166, n_542);
  not gc166 (wc166, n_543);
  or g1944 (n_1854, n_601, wc167);
  not gc167 (wc167, n_605);
  or g1945 (n_1855, wc168, n_597);
  not gc168 (wc168, n_598);
  and g1946 (n_1856, wc169, n_500);
  not gc169 (wc169, B[6]);
  and g1947 (n_1857, n_317, n_548);
  and g1948 (n_1858, n_460, n_603);
  or g1949 (n_1859, n_1841, wc170);
  not gc170 (wc170, n_512);
  or g1950 (n_1860, n_570, wc171);
  not gc171 (wc171, n_563);
  or g1951 (n_1861, n_625, wc172);
  not gc172 (wc172, n_618);
  or g1952 (n_487, wc173, n_1856);
  not gc173 (wc173, n_1859);
  or g1953 (n_535, wc174, n_1857);
  not gc174 (wc174, n_1860);
  or g1954 (n_1862, wc175, n_1858);
  not gc175 (wc175, n_1861);
  or g1955 (n_81, wc176, n_1831);
  not gc176 (wc176, n_1862);
  and g1956 (n_80, wc177, n_487);
  not gc177 (wc177, n_535);
  or g1957 (QUOTIENT[11], wc178, n_535);
  not gc178 (wc178, n_81);
  or g1958 (QUOTIENT[10], n_80, wc179);
  not gc179 (wc179, n_81);
  or g1959 (n_89, wc180, wc182, wc183, wc184);
  and gc185 (wc184, wc185, n_77);
  not gc184 (wc185, n_81);
  and gc183 (wc183, n_76, n_82);
  and gc182 (wc182, n_80, n_75);
  and gc181 (wc180, wc181, n_65);
  not gc180 (wc181, n_487);
  or g1960 (n_87, wc186, wc188, wc189, wc190);
  and gc191 (wc190, wc191, n_71);
  not gc190 (wc191, n_81);
  and gc189 (wc189, n_70, n_82);
  and gc188 (wc188, n_80, n_69);
  and gc187 (wc186, wc187, n_63);
  not gc186 (wc187, n_487);
  or g1961 (n_88, wc192, wc194, wc195, wc196);
  and gc197 (wc196, wc197, n_74);
  not gc196 (wc197, n_81);
  and gc195 (wc195, n_73, n_82);
  and gc194 (wc194, n_80, n_72);
  and gc193 (wc192, wc193, n_64);
  not gc192 (wc193, n_487);
  or g1962 (n_85, wc198, wc200, wc202, wc203);
  and gc205 (wc203, wc204, wc205);
  not gc204 (wc205, n_1764);
  not gc203 (wc204, n_81);
  and gc202 (wc202, A[10], n_82);
  and gc201 (wc200, n_80, wc201);
  not gc200 (wc201, n_1764);
  and gc199 (wc198, A[10], wc199);
  not gc198 (wc199, n_487);
  or g1963 (n_86, wc206, wc208, wc209, wc210);
  and gc211 (wc210, wc211, n_68);
  not gc210 (wc211, n_81);
  and gc209 (wc209, n_1800, n_82);
  and gc208 (wc208, n_80, n_67);
  and gc207 (wc206, A[11], wc207);
  not gc206 (wc207, n_487);
  and g1964 (n_674, B[6], wc212);
  not gc212 (wc212, n_89);
  or g1965 (n_662, B[4], wc213);
  not gc213 (wc213, n_87);
  and g1966 (n_663, B[5], wc214);
  not gc214 (wc214, n_88);
  or g1967 (n_664, B[5], wc215);
  not gc215 (wc215, n_88);
  or g1968 (n_676, B[6], wc216);
  not gc216 (wc216, n_89);
  or g1969 (n_656, B[2], wc217);
  not gc217 (wc217, n_85);
  and g1970 (n_657, B[3], wc218);
  not gc218 (wc218, n_86);
  or g1971 (n_658, B[3], wc219);
  not gc219 (wc219, n_86);
  and g1972 (n_661, B[2], wc220);
  not gc220 (wc220, n_85);
  and g1973 (n_667, B[4], wc221);
  not gc221 (wc221, n_87);
  or g1974 (n_721, B[3], wc222);
  not gc222 (wc222, n_87);
  and g1975 (n_722, B[4], wc223);
  not gc223 (wc223, n_88);
  or g1976 (n_723, B[4], wc224);
  not gc224 (wc224, n_88);
  and g1977 (n_729, B[5], wc225);
  not gc225 (wc225, n_89);
  or g1978 (n_727, B[5], wc226);
  not gc226 (wc226, n_89);
  or g1979 (n_715, B[1], wc227);
  not gc227 (wc227, n_85);
  and g1980 (n_716, B[2], wc228);
  not gc228 (wc228, n_86);
  or g1981 (n_717, B[2], wc229);
  not gc229 (wc229, n_86);
  and g1982 (n_720, B[1], wc230);
  not gc230 (wc230, n_85);
  and g1983 (n_726, B[3], wc231);
  not gc231 (wc231, n_87);
  or g1984 (n_788, wc232, n_43);
  not gc232 (wc232, n_87);
  and g1985 (n_789, wc233, n_44);
  not gc233 (wc233, n_88);
  or g1986 (n_790, wc234, n_44);
  not gc234 (wc234, n_88);
  and g1987 (n_796, wc235, n_45);
  not gc235 (wc235, n_89);
  or g1988 (n_794, wc236, n_45);
  not gc236 (wc236, n_89);
  or g1989 (n_782, wc237, n_1794);
  not gc237 (wc237, n_85);
  and g1990 (n_783, wc238, n_42);
  not gc238 (wc238, n_86);
  or g1991 (n_784, wc239, n_42);
  not gc239 (wc239, n_86);
  and g1992 (n_787, wc240, n_1794);
  not gc240 (wc240, n_85);
  and g1993 (n_793, wc241, n_43);
  not gc241 (wc241, n_87);
  and g1994 (n_675, n_664, wc242);
  not gc242 (wc242, n_665);
  and g1995 (n_1865, n_658, wc243);
  not gc243 (wc243, n_659);
  or g1996 (n_1866, n_674, wc244);
  not gc244 (wc244, n_679);
  and g1997 (n_736, n_723, wc245);
  not gc245 (wc245, n_724);
  and g1998 (n_1867, n_717, wc246);
  not gc246 (wc246, n_718);
  and g1999 (n_803, n_790, wc247);
  not gc247 (wc247, n_791);
  and g2000 (n_1868, n_784, wc248);
  not gc248 (wc248, n_785);
  or g2001 (n_1869, wc249, n_674);
  not gc249 (wc249, n_676);
  or g2002 (n_1870, wc250, n_729);
  not gc250 (wc250, n_727);
  or g2003 (n_1871, wc251, n_796);
  not gc251 (wc251, n_794);
  or g2004 (n_1872, n_661, wc252);
  not gc252 (wc252, n_656);
  or g2005 (n_1873, n_720, wc253);
  not gc253 (wc253, n_715);
  or g2006 (n_1874, n_787, wc254);
  not gc254 (wc254, n_782);
  or g2007 (n_1875, n_661, wc255);
  not gc255 (wc255, n_668);
  or g2008 (n_1876, wc256, n_657);
  not gc256 (wc256, n_658);
  or g2009 (n_1877, n_720, wc257);
  not gc257 (wc257, n_730);
  or g2010 (n_1878, wc258, n_716);
  not gc258 (wc258, n_717);
  or g2011 (n_1879, n_787, wc259);
  not gc259 (wc259, n_797);
  or g2012 (n_1880, wc260, n_783);
  not gc260 (wc260, n_784);
  or g2013 (n_1881, n_667, wc261);
  not gc261 (wc261, n_662);
  or g2014 (n_1882, n_726, wc262);
  not gc262 (wc262, n_721);
  or g2015 (n_1883, n_793, wc263);
  not gc263 (wc263, n_788);
  or g2016 (n_1884, wc264, n_663);
  not gc264 (wc264, n_664);
  or g2017 (n_1885, wc265, n_722);
  not gc265 (wc265, n_723);
  or g2018 (n_1886, wc266, n_789);
  not gc266 (wc266, n_790);
  and g2019 (n_1887, wc267, n_741);
  not gc267 (wc267, n_736);
  and g2020 (n_1888, wc268, n_808);
  not gc268 (wc268, n_803);
  and g2021 (n_1889, n_676, wc269);
  not gc269 (wc269, n_677);
  or g2022 (n_1890, n_1866, wc270);
  not gc270 (wc270, n_681);
  or g2023 (n_1891, n_752, wc271);
  not gc271 (wc271, n_744);
  or g2024 (n_1892, n_819, wc272);
  not gc272 (wc272, n_811);
  or g2025 (n_1893, n_667, wc273);
  not gc273 (wc273, n_681);
  or g2026 (n_1894, n_726, wc274);
  not gc274 (wc274, n_744);
  or g2027 (n_1895, n_793, wc275);
  not gc275 (wc275, n_811);
  or g2028 (n_111, n_1831, wc276);
  not gc276 (wc276, n_823);
  and g2029 (n_110, wc277, n_650);
  not gc277 (wc277, n_709);
  or g2030 (QUOTIENT[9], wc278, n_709);
  not gc278 (wc278, n_111);
  or g2031 (QUOTIENT[8], n_110, wc279);
  not gc279 (wc279, n_111);
  or g2032 (n_121, wc280, wc282, wc283, wc284);
  and gc285 (wc284, wc285, n_107);
  not gc284 (wc285, n_111);
  and gc283 (wc283, n_106, n_112);
  and gc282 (wc282, n_110, n_105);
  and gc281 (wc280, n_89, wc281);
  not gc280 (wc281, n_650);
  or g2033 (n_117, wc286, wc288, wc289, wc290);
  and gc291 (wc290, wc291, n_95);
  not gc290 (wc291, n_111);
  and gc289 (wc289, n_94, n_112);
  and gc288 (wc288, n_110, n_93);
  and gc287 (wc286, n_85, wc287);
  not gc286 (wc287, n_650);
  or g2034 (n_118, wc292, wc294, wc295, wc296);
  and gc297 (wc296, wc297, n_98);
  not gc296 (wc297, n_111);
  and gc295 (wc295, n_97, n_112);
  and gc294 (wc294, n_110, n_96);
  and gc293 (wc292, n_86, wc293);
  not gc292 (wc293, n_650);
  or g2035 (n_119, wc298, wc300, wc301, wc302);
  and gc303 (wc302, wc303, n_101);
  not gc302 (wc303, n_111);
  and gc301 (wc301, n_100, n_112);
  and gc300 (wc300, n_110, n_99);
  and gc299 (wc298, n_87, wc299);
  not gc298 (wc299, n_650);
  or g2036 (n_120, wc304, wc306, wc307, wc308);
  and gc309 (wc308, wc309, n_104);
  not gc308 (wc309, n_111);
  and gc307 (wc307, n_103, n_112);
  and gc306 (wc306, n_110, n_102);
  and gc305 (wc304, n_88, wc305);
  not gc304 (wc305, n_650);
  or g2037 (n_115, wc310, wc312, wc314, wc315);
  and gc317 (wc315, wc316, wc317);
  not gc316 (wc317, n_1766);
  not gc315 (wc316, n_111);
  and gc314 (wc314, A[8], n_112);
  and gc313 (wc312, n_110, wc313);
  not gc312 (wc313, n_1766);
  and gc311 (wc310, A[8], wc311);
  not gc310 (wc311, n_650);
  or g2038 (n_116, wc318, wc320, wc321, wc322);
  and gc323 (wc322, wc323, n_92);
  not gc322 (wc323, n_111);
  and gc321 (wc321, n_1803, n_112);
  and gc320 (wc320, n_110, n_91);
  and gc319 (wc318, A[9], wc319);
  not gc318 (wc319, n_650);
  or g2039 (n_858, B[4], wc324);
  not gc324 (wc324, n_117);
  and g2040 (n_859, B[5], wc325);
  not gc325 (wc325, n_118);
  or g2041 (n_860, B[5], wc326);
  not gc326 (wc326, n_118);
  and g2042 (n_865, B[6], wc327);
  not gc327 (wc327, n_119);
  or g2043 (n_864, B[6], wc328);
  not gc328 (wc328, n_119);
  or g2044 (n_852, B[2], wc329);
  not gc329 (wc329, n_115);
  and g2045 (n_853, B[3], wc330);
  not gc330 (wc330, n_116);
  or g2046 (n_854, B[3], wc331);
  not gc331 (wc331, n_116);
  and g2047 (n_857, B[2], wc332);
  not gc332 (wc332, n_115);
  and g2048 (n_863, B[4], wc333);
  not gc333 (wc333, n_117);
  or g2049 (n_926, B[3], wc334);
  not gc334 (wc334, n_117);
  and g2050 (n_927, B[4], wc335);
  not gc335 (wc335, n_118);
  or g2051 (n_928, B[4], wc336);
  not gc336 (wc336, n_118);
  and g2052 (n_937, B[5], wc337);
  not gc337 (wc337, n_119);
  and g2053 (n_933, B[6], wc338);
  not gc338 (wc338, n_120);
  or g2054 (n_932, B[5], wc339);
  not gc339 (wc339, n_119);
  or g2055 (n_1898, B[6], wc340);
  not gc340 (wc340, n_120);
  or g2056 (n_920, B[1], wc341);
  not gc341 (wc341, n_115);
  and g2057 (n_921, B[2], wc342);
  not gc342 (wc342, n_116);
  or g2058 (n_922, B[2], wc343);
  not gc343 (wc343, n_116);
  and g2059 (n_925, B[1], wc344);
  not gc344 (wc344, n_115);
  and g2060 (n_931, B[3], wc345);
  not gc345 (wc345, n_117);
  or g2061 (n_1899, wc346, n_1831);
  not gc346 (wc346, n_121);
  or g2062 (n_1006, wc347, n_43);
  not gc347 (wc347, n_117);
  and g2063 (n_1007, wc348, n_44);
  not gc348 (wc348, n_118);
  or g2064 (n_1008, wc349, n_44);
  not gc349 (wc349, n_118);
  and g2065 (n_1017, wc350, n_45);
  not gc350 (wc350, n_119);
  and g2066 (n_1013, wc351, n_46);
  not gc351 (wc351, n_120);
  or g2067 (n_1012, wc352, n_45);
  not gc352 (wc352, n_119);
  or g2068 (n_1900, wc353, n_46);
  not gc353 (wc353, n_120);
  or g2069 (n_1000, wc354, n_1794);
  not gc354 (wc354, n_115);
  and g2070 (n_1001, wc355, n_42);
  not gc355 (wc355, n_116);
  or g2071 (n_1002, wc356, n_42);
  not gc356 (wc356, n_116);
  and g2072 (n_1005, wc357, n_1794);
  not gc357 (wc357, n_115);
  and g2073 (n_1011, wc358, n_43);
  not gc358 (wc358, n_117);
  and g2074 (n_1901, wc359, n_1831);
  not gc359 (wc359, n_121);
  and g2075 (n_872, n_860, wc360);
  not gc360 (wc360, n_861);
  and g2076 (n_1902, n_864, wc361);
  not gc361 (wc361, n_120);
  and g2077 (n_1903, n_854, wc362);
  not gc362 (wc362, n_855);
  or g2078 (n_1904, n_865, wc363);
  not gc363 (wc363, n_875);
  and g2079 (n_944, n_928, wc364);
  not gc364 (wc364, n_929);
  and g2080 (n_1905, n_1898, wc365);
  not gc365 (wc365, n_935);
  and g2081 (n_1906, n_922, wc366);
  not gc366 (wc366, n_923);
  and g2082 (n_1024, n_1008, wc367);
  not gc367 (wc367, n_1009);
  and g2083 (n_1907, n_1900, wc368);
  not gc368 (wc368, n_1015);
  and g2084 (n_1908, n_1002, wc369);
  not gc369 (wc369, n_1003);
  or g2085 (n_1909, wc370, n_865);
  not gc370 (wc370, n_864);
  or g2086 (n_1910, wc371, n_937);
  not gc371 (wc371, n_932);
  or g2087 (n_1911, wc372, n_1017);
  not gc372 (wc372, n_1012);
  or g2088 (n_1912, n_857, wc373);
  not gc373 (wc373, n_852);
  or g2089 (n_1913, n_925, wc374);
  not gc374 (wc374, n_920);
  or g2090 (n_1914, n_1005, wc375);
  not gc375 (wc375, n_1000);
  or g2091 (n_1915, n_857, wc376);
  not gc376 (wc376, n_866);
  or g2092 (n_1916, wc377, n_853);
  not gc377 (wc377, n_854);
  or g2093 (n_1917, n_925, wc378);
  not gc378 (wc378, n_938);
  or g2094 (n_1918, wc379, n_921);
  not gc379 (wc379, n_922);
  or g2095 (n_1919, n_1005, wc380);
  not gc380 (wc380, n_1018);
  or g2096 (n_1920, wc381, n_1001);
  not gc381 (wc381, n_1002);
  or g2097 (n_1921, n_863, wc382);
  not gc382 (wc382, n_858);
  or g2098 (n_1922, n_931, wc383);
  not gc383 (wc383, n_926);
  or g2099 (n_1923, n_1011, wc384);
  not gc384 (wc384, n_1006);
  or g2100 (n_1924, wc385, n_859);
  not gc385 (wc385, n_860);
  or g2101 (n_1925, wc386, n_927);
  not gc386 (wc386, n_928);
  or g2102 (n_1926, wc387, n_1007);
  not gc387 (wc387, n_1008);
  and g2103 (n_1927, wc388, n_949);
  not gc388 (wc388, n_944);
  and g2104 (n_1928, wc389, n_1029);
  not gc389 (wc389, n_1024);
  and g2105 (n_1929, n_1902, wc390);
  not gc390 (wc390, n_878);
  or g2106 (n_1930, n_1904, wc391);
  not gc391 (wc391, n_880);
  and g2107 (n_1931, wc392, n_1905);
  not gc392 (wc392, n_1927);
  or g2108 (n_1932, n_962, wc393);
  not gc393 (wc393, n_954);
  and g2109 (n_1933, wc394, n_1907);
  not gc394 (wc394, n_1928);
  or g2110 (n_1934, n_1042, wc395);
  not gc395 (wc395, n_1034);
  or g2111 (n_1935, n_863, wc396);
  not gc396 (wc396, n_880);
  or g2112 (n_1936, n_931, wc397);
  not gc397 (wc397, n_954);
  or g2113 (n_1937, n_1011, wc398);
  not gc398 (wc398, n_1034);
  or g2114 (n_1938, n_1901, wc399);
  not gc399 (wc399, n_1047);
  or g2115 (n_846, n_889, n_121);
  or g2116 (n_914, n_966, n_121);
  and g2117 (n_147, wc400, n_846);
  not gc400 (wc400, n_914);
  and g2118 (n_150, n_914, wc401);
  not gc401 (wc401, n_151);
  or g2119 (QUOTIENT[7], n_151, n_914);
  or g2120 (n_161, wc402, wc404, wc405, wc406);
  and gc406 (wc406, n_139, n_151);
  and gc405 (wc405, n_150, n_138);
  and gc404 (wc404, n_147, n_137);
  and gc403 (wc402, wc403, n_119);
  not gc402 (wc403, n_846);
  or g2121 (n_157, wc407, wc409, wc410, wc411);
  and gc411 (wc411, n_127, n_151);
  and gc410 (wc410, n_150, n_126);
  and gc409 (wc409, n_147, n_125);
  and gc408 (wc407, wc408, n_115);
  not gc407 (wc408, n_846);
  or g2122 (n_158, wc412, wc414, wc415, wc416);
  and gc416 (wc416, n_130, n_151);
  and gc415 (wc415, n_150, n_129);
  and gc414 (wc414, n_147, n_128);
  and gc413 (wc412, wc413, n_116);
  not gc412 (wc413, n_846);
  or g2123 (n_159, wc417, wc419, wc420, wc421);
  and gc421 (wc421, n_133, n_151);
  and gc420 (wc420, n_150, n_132);
  and gc419 (wc419, n_147, n_131);
  and gc418 (wc417, wc418, n_117);
  not gc417 (wc418, n_846);
  or g2124 (n_160, wc422, wc424, wc425, wc426);
  and gc426 (wc426, n_136, n_151);
  and gc425 (wc425, n_150, n_135);
  and gc424 (wc424, n_147, n_134);
  and gc423 (wc422, wc423, n_118);
  not gc422 (wc423, n_846);
  or g2125 (n_155, wc427, wc429, wc431, wc432);
  and gc433 (wc432, wc433, n_151);
  not gc432 (wc433, n_1768);
  and gc431 (wc431, A[6], n_150);
  and gc430 (wc429, n_147, wc430);
  not gc429 (wc430, n_1768);
  and gc428 (wc427, A[6], wc428);
  not gc427 (wc428, n_846);
  or g2126 (n_156, wc434, wc436, wc437, wc438);
  and gc438 (wc438, n_124, n_151);
  and gc437 (wc437, n_150, n_1806);
  and gc436 (wc436, n_147, n_123);
  and gc435 (wc434, A[7], wc435);
  not gc434 (wc435, n_846);
  or g2127 (n_1087, B[4], wc439);
  not gc439 (wc439, n_157);
  and g2128 (n_1088, B[5], wc440);
  not gc440 (wc440, n_158);
  or g2129 (n_1089, B[5], wc441);
  not gc441 (wc441, n_158);
  and g2130 (n_1094, B[6], wc442);
  not gc442 (wc442, n_159);
  or g2131 (n_1093, B[6], wc443);
  not gc443 (wc443, n_159);
  or g2132 (n_1081, B[2], wc444);
  not gc444 (wc444, n_155);
  and g2133 (n_1082, B[3], wc445);
  not gc445 (wc445, n_156);
  or g2134 (n_1083, B[3], wc446);
  not gc446 (wc446, n_156);
  and g2135 (n_1086, B[2], wc447);
  not gc447 (wc447, n_155);
  and g2136 (n_1092, B[4], wc448);
  not gc448 (wc448, n_157);
  or g2137 (n_1155, B[3], wc449);
  not gc449 (wc449, n_157);
  and g2138 (n_1156, B[4], wc450);
  not gc450 (wc450, n_158);
  or g2139 (n_1157, B[4], wc451);
  not gc451 (wc451, n_158);
  and g2140 (n_1166, B[5], wc452);
  not gc452 (wc452, n_159);
  and g2141 (n_1162, B[6], wc453);
  not gc453 (wc453, n_160);
  or g2142 (n_1161, B[5], wc454);
  not gc454 (wc454, n_159);
  or g2143 (n_1940, B[6], wc455);
  not gc455 (wc455, n_160);
  or g2144 (n_1149, B[1], wc456);
  not gc456 (wc456, n_155);
  and g2145 (n_1150, B[2], wc457);
  not gc457 (wc457, n_156);
  or g2146 (n_1151, B[2], wc458);
  not gc458 (wc458, n_156);
  and g2147 (n_1154, B[1], wc459);
  not gc459 (wc459, n_155);
  and g2148 (n_1160, B[3], wc460);
  not gc460 (wc460, n_157);
  or g2149 (n_1941, wc461, n_1831);
  not gc461 (wc461, n_161);
  or g2150 (n_1235, wc462, n_43);
  not gc462 (wc462, n_157);
  and g2151 (n_1236, wc463, n_44);
  not gc463 (wc463, n_158);
  or g2152 (n_1237, wc464, n_44);
  not gc464 (wc464, n_158);
  and g2153 (n_1246, wc465, n_45);
  not gc465 (wc465, n_159);
  and g2154 (n_1242, wc466, n_46);
  not gc466 (wc466, n_160);
  or g2155 (n_1241, wc467, n_45);
  not gc467 (wc467, n_159);
  or g2156 (n_1942, wc468, n_46);
  not gc468 (wc468, n_160);
  or g2157 (n_1229, wc469, n_1794);
  not gc469 (wc469, n_155);
  and g2158 (n_1230, wc470, n_42);
  not gc470 (wc470, n_156);
  or g2159 (n_1231, wc471, n_42);
  not gc471 (wc471, n_156);
  and g2160 (n_1234, wc472, n_1794);
  not gc472 (wc472, n_155);
  and g2161 (n_1240, wc473, n_43);
  not gc473 (wc473, n_157);
  and g2162 (n_1943, wc474, n_1831);
  not gc474 (wc474, n_161);
  and g2163 (n_1101, n_1089, wc475);
  not gc475 (wc475, n_1090);
  and g2164 (n_1944, n_1093, wc476);
  not gc476 (wc476, n_160);
  and g2165 (n_1945, n_1083, wc477);
  not gc477 (wc477, n_1084);
  or g2166 (n_1946, n_1094, wc478);
  not gc478 (wc478, n_1104);
  and g2167 (n_1173, n_1157, wc479);
  not gc479 (wc479, n_1158);
  and g2168 (n_1947, n_1940, wc480);
  not gc480 (wc480, n_1164);
  and g2169 (n_1948, n_1151, wc481);
  not gc481 (wc481, n_1152);
  and g2170 (n_1253, n_1237, wc482);
  not gc482 (wc482, n_1238);
  and g2171 (n_1949, n_1942, wc483);
  not gc483 (wc483, n_1244);
  and g2172 (n_1950, n_1231, wc484);
  not gc484 (wc484, n_1232);
  or g2173 (n_1951, wc485, n_1094);
  not gc485 (wc485, n_1093);
  or g2174 (n_1952, wc486, n_1166);
  not gc486 (wc486, n_1161);
  or g2175 (n_1953, wc487, n_1246);
  not gc487 (wc487, n_1241);
  or g2176 (n_1954, n_1086, wc488);
  not gc488 (wc488, n_1081);
  or g2177 (n_1955, n_1154, wc489);
  not gc489 (wc489, n_1149);
  or g2178 (n_1956, n_1234, wc490);
  not gc490 (wc490, n_1229);
  or g2179 (n_1957, n_1086, wc491);
  not gc491 (wc491, n_1095);
  or g2180 (n_1958, wc492, n_1082);
  not gc492 (wc492, n_1083);
  or g2181 (n_1959, n_1154, wc493);
  not gc493 (wc493, n_1167);
  or g2182 (n_1960, wc494, n_1150);
  not gc494 (wc494, n_1151);
  or g2183 (n_1961, n_1234, wc495);
  not gc495 (wc495, n_1247);
  or g2184 (n_1962, wc496, n_1230);
  not gc496 (wc496, n_1231);
  or g2185 (n_1963, n_1092, wc497);
  not gc497 (wc497, n_1087);
  or g2186 (n_1964, n_1160, wc498);
  not gc498 (wc498, n_1155);
  or g2187 (n_1965, n_1240, wc499);
  not gc499 (wc499, n_1235);
  or g2188 (n_1966, wc500, n_1088);
  not gc500 (wc500, n_1089);
  or g2189 (n_1967, wc501, n_1156);
  not gc501 (wc501, n_1157);
  or g2190 (n_1968, wc502, n_1236);
  not gc502 (wc502, n_1237);
  and g2191 (n_1969, wc503, n_1178);
  not gc503 (wc503, n_1173);
  and g2192 (n_1970, wc504, n_1258);
  not gc504 (wc504, n_1253);
  and g2193 (n_1971, n_1944, wc505);
  not gc505 (wc505, n_1107);
  or g2194 (n_1972, n_1946, wc506);
  not gc506 (wc506, n_1109);
  and g2195 (n_1973, wc507, n_1947);
  not gc507 (wc507, n_1969);
  or g2196 (n_1974, n_1191, wc508);
  not gc508 (wc508, n_1183);
  and g2197 (n_1975, wc509, n_1949);
  not gc509 (wc509, n_1970);
  or g2198 (n_1976, n_1271, wc510);
  not gc510 (wc510, n_1263);
  or g2199 (n_1977, n_1092, wc511);
  not gc511 (wc511, n_1109);
  or g2200 (n_1978, n_1160, wc512);
  not gc512 (wc512, n_1183);
  or g2201 (n_1979, n_1240, wc513);
  not gc513 (wc513, n_1263);
  or g2202 (n_1980, n_1943, wc514);
  not gc514 (wc514, n_1276);
  or g2203 (n_1075, n_1118, n_161);
  or g2204 (n_1143, n_1195, n_161);
  and g2205 (n_192, wc515, n_1075);
  not gc515 (wc515, n_1143);
  and g2206 (n_195, n_1143, wc516);
  not gc516 (wc516, n_196);
  or g2207 (QUOTIENT[5], n_196, n_1143);
  or g2208 (n_206, wc517, wc519, wc520, wc521);
  and gc521 (wc521, n_182, n_196);
  and gc520 (wc520, n_195, n_181);
  and gc519 (wc519, n_192, n_180);
  and gc518 (wc517, wc518, n_159);
  not gc517 (wc518, n_1075);
  or g2209 (n_202, wc522, wc524, wc525, wc526);
  and gc526 (wc526, n_170, n_196);
  and gc525 (wc525, n_195, n_169);
  and gc524 (wc524, n_192, n_168);
  and gc523 (wc522, wc523, n_155);
  not gc522 (wc523, n_1075);
  or g2210 (n_203, wc527, wc529, wc530, wc531);
  and gc531 (wc531, n_173, n_196);
  and gc530 (wc530, n_195, n_172);
  and gc529 (wc529, n_192, n_171);
  and gc528 (wc527, wc528, n_156);
  not gc527 (wc528, n_1075);
  or g2211 (n_204, wc532, wc534, wc535, wc536);
  and gc536 (wc536, n_176, n_196);
  and gc535 (wc535, n_195, n_175);
  and gc534 (wc534, n_192, n_174);
  and gc533 (wc532, wc533, n_157);
  not gc532 (wc533, n_1075);
  or g2212 (n_205, wc537, wc539, wc540, wc541);
  and gc541 (wc541, n_179, n_196);
  and gc540 (wc540, n_195, n_178);
  and gc539 (wc539, n_192, n_177);
  and gc538 (wc537, wc538, n_158);
  not gc537 (wc538, n_1075);
  or g2213 (n_200, wc542, wc544, wc546, wc547);
  and gc548 (wc547, wc548, n_196);
  not gc547 (wc548, n_1770);
  and gc546 (wc546, A[4], n_195);
  and gc545 (wc544, n_192, wc545);
  not gc544 (wc545, n_1770);
  and gc543 (wc542, A[4], wc543);
  not gc542 (wc543, n_1075);
  or g2214 (n_201, wc549, wc551, wc552, wc553);
  and gc553 (wc553, n_167, n_196);
  and gc552 (wc552, n_195, n_1809);
  and gc551 (wc551, n_192, n_165);
  and gc550 (wc549, A[5], wc550);
  not gc549 (wc550, n_1075);
  or g2215 (n_1316, B[4], wc554);
  not gc554 (wc554, n_202);
  and g2216 (n_1317, B[5], wc555);
  not gc555 (wc555, n_203);
  or g2217 (n_1318, B[5], wc556);
  not gc556 (wc556, n_203);
  and g2218 (n_1323, B[6], wc557);
  not gc557 (wc557, n_204);
  or g2219 (n_1322, B[6], wc558);
  not gc558 (wc558, n_204);
  or g2220 (n_1310, B[2], wc559);
  not gc559 (wc559, n_200);
  and g2221 (n_1311, B[3], wc560);
  not gc560 (wc560, n_201);
  or g2222 (n_1312, B[3], wc561);
  not gc561 (wc561, n_201);
  and g2223 (n_1315, B[2], wc562);
  not gc562 (wc562, n_200);
  and g2224 (n_1321, B[4], wc563);
  not gc563 (wc563, n_202);
  or g2225 (n_1384, B[3], wc564);
  not gc564 (wc564, n_202);
  and g2226 (n_1385, B[4], wc565);
  not gc565 (wc565, n_203);
  or g2227 (n_1386, B[4], wc566);
  not gc566 (wc566, n_203);
  and g2228 (n_1395, B[5], wc567);
  not gc567 (wc567, n_204);
  and g2229 (n_1391, B[6], wc568);
  not gc568 (wc568, n_205);
  or g2230 (n_1390, B[5], wc569);
  not gc569 (wc569, n_204);
  or g2231 (n_1982, B[6], wc570);
  not gc570 (wc570, n_205);
  or g2232 (n_1378, B[1], wc571);
  not gc571 (wc571, n_200);
  and g2233 (n_1379, B[2], wc572);
  not gc572 (wc572, n_201);
  or g2234 (n_1380, B[2], wc573);
  not gc573 (wc573, n_201);
  and g2235 (n_1383, B[1], wc574);
  not gc574 (wc574, n_200);
  and g2236 (n_1389, B[3], wc575);
  not gc575 (wc575, n_202);
  or g2237 (n_1983, wc576, n_1831);
  not gc576 (wc576, n_206);
  or g2238 (n_1464, wc577, n_43);
  not gc577 (wc577, n_202);
  and g2239 (n_1465, wc578, n_44);
  not gc578 (wc578, n_203);
  or g2240 (n_1466, wc579, n_44);
  not gc579 (wc579, n_203);
  and g2241 (n_1475, wc580, n_45);
  not gc580 (wc580, n_204);
  and g2242 (n_1471, wc581, n_46);
  not gc581 (wc581, n_205);
  or g2243 (n_1470, wc582, n_45);
  not gc582 (wc582, n_204);
  or g2244 (n_1984, wc583, n_46);
  not gc583 (wc583, n_205);
  or g2245 (n_1458, wc584, n_1794);
  not gc584 (wc584, n_200);
  and g2246 (n_1459, wc585, n_42);
  not gc585 (wc585, n_201);
  or g2247 (n_1460, wc586, n_42);
  not gc586 (wc586, n_201);
  and g2248 (n_1463, wc587, n_1794);
  not gc587 (wc587, n_200);
  and g2249 (n_1469, wc588, n_43);
  not gc588 (wc588, n_202);
  and g2250 (n_1985, wc589, n_1831);
  not gc589 (wc589, n_206);
  and g2251 (n_1330, n_1318, wc590);
  not gc590 (wc590, n_1319);
  and g2252 (n_1986, n_1322, wc591);
  not gc591 (wc591, n_205);
  and g2253 (n_1987, n_1312, wc592);
  not gc592 (wc592, n_1313);
  or g2254 (n_1988, n_1323, wc593);
  not gc593 (wc593, n_1333);
  and g2255 (n_1402, n_1386, wc594);
  not gc594 (wc594, n_1387);
  and g2256 (n_1989, n_1982, wc595);
  not gc595 (wc595, n_1393);
  and g2257 (n_1990, n_1380, wc596);
  not gc596 (wc596, n_1381);
  and g2258 (n_1482, n_1466, wc597);
  not gc597 (wc597, n_1467);
  and g2259 (n_1991, n_1984, wc598);
  not gc598 (wc598, n_1473);
  and g2260 (n_1992, n_1460, wc599);
  not gc599 (wc599, n_1461);
  or g2261 (n_1993, wc600, n_1323);
  not gc600 (wc600, n_1322);
  or g2262 (n_1994, wc601, n_1395);
  not gc601 (wc601, n_1390);
  or g2263 (n_1995, wc602, n_1475);
  not gc602 (wc602, n_1470);
  or g2264 (n_1996, n_1315, wc603);
  not gc603 (wc603, n_1310);
  or g2265 (n_1997, n_1383, wc604);
  not gc604 (wc604, n_1378);
  or g2266 (n_1998, n_1463, wc605);
  not gc605 (wc605, n_1458);
  or g2267 (n_1999, n_1315, wc606);
  not gc606 (wc606, n_1324);
  or g2268 (n_2000, wc607, n_1311);
  not gc607 (wc607, n_1312);
  or g2269 (n_2001, n_1383, wc608);
  not gc608 (wc608, n_1396);
  or g2270 (n_2002, wc609, n_1379);
  not gc609 (wc609, n_1380);
  or g2271 (n_2003, n_1463, wc610);
  not gc610 (wc610, n_1476);
  or g2272 (n_2004, wc611, n_1459);
  not gc611 (wc611, n_1460);
  or g2273 (n_2005, n_1321, wc612);
  not gc612 (wc612, n_1316);
  or g2274 (n_2006, n_1389, wc613);
  not gc613 (wc613, n_1384);
  or g2275 (n_2007, n_1469, wc614);
  not gc614 (wc614, n_1464);
  or g2276 (n_2008, wc615, n_1317);
  not gc615 (wc615, n_1318);
  or g2277 (n_2009, wc616, n_1385);
  not gc616 (wc616, n_1386);
  or g2278 (n_2010, wc617, n_1465);
  not gc617 (wc617, n_1466);
  and g2279 (n_2011, wc618, n_1407);
  not gc618 (wc618, n_1402);
  and g2280 (n_2012, wc619, n_1487);
  not gc619 (wc619, n_1482);
  and g2281 (n_2013, n_1986, wc620);
  not gc620 (wc620, n_1336);
  or g2282 (n_2014, n_1988, wc621);
  not gc621 (wc621, n_1338);
  and g2283 (n_2015, wc622, n_1989);
  not gc622 (wc622, n_2011);
  or g2284 (n_2016, n_1420, wc623);
  not gc623 (wc623, n_1412);
  and g2285 (n_2017, wc624, n_1991);
  not gc624 (wc624, n_2012);
  or g2286 (n_2018, n_1500, wc625);
  not gc625 (wc625, n_1492);
  or g2287 (n_2019, n_1321, wc626);
  not gc626 (wc626, n_1338);
  or g2288 (n_2020, n_1389, wc627);
  not gc627 (wc627, n_1412);
  or g2289 (n_2021, n_1469, wc628);
  not gc628 (wc628, n_1492);
  or g2290 (n_2022, n_1985, wc629);
  not gc629 (wc629, n_1505);
  or g2291 (n_1304, n_1347, n_206);
  or g2292 (n_1372, n_1424, n_206);
  and g2293 (n_237, wc630, n_1304);
  not gc630 (wc630, n_1372);
  and g2294 (n_240, n_1372, wc631);
  not gc631 (wc631, n_241);
  or g2295 (QUOTIENT[3], n_241, n_1372);
  or g2296 (n_251, wc632, wc634, wc635, wc636);
  and gc636 (wc636, n_227, n_241);
  and gc635 (wc635, n_240, n_226);
  and gc634 (wc634, n_237, n_225);
  and gc633 (wc632, wc633, n_204);
  not gc632 (wc633, n_1304);
  or g2297 (n_247, wc637, wc639, wc640, wc641);
  and gc641 (wc641, n_215, n_241);
  and gc640 (wc640, n_240, n_214);
  and gc639 (wc639, n_237, n_213);
  and gc638 (wc637, wc638, n_200);
  not gc637 (wc638, n_1304);
  or g2298 (n_248, wc642, wc644, wc645, wc646);
  and gc646 (wc646, n_218, n_241);
  and gc645 (wc645, n_240, n_217);
  and gc644 (wc644, n_237, n_216);
  and gc643 (wc642, wc643, n_201);
  not gc642 (wc643, n_1304);
  or g2299 (n_249, wc647, wc649, wc650, wc651);
  and gc651 (wc651, n_221, n_241);
  and gc650 (wc650, n_240, n_220);
  and gc649 (wc649, n_237, n_219);
  and gc648 (wc647, wc648, n_202);
  not gc647 (wc648, n_1304);
  or g2300 (n_250, wc652, wc654, wc655, wc656);
  and gc656 (wc656, n_224, n_241);
  and gc655 (wc655, n_240, n_223);
  and gc654 (wc654, n_237, n_222);
  and gc653 (wc652, wc653, n_203);
  not gc652 (wc653, n_1304);
  or g2301 (n_245, wc657, wc659, wc661, wc662);
  and gc663 (wc662, wc663, n_241);
  not gc662 (wc663, n_1772);
  and gc661 (wc661, A[2], n_240);
  and gc660 (wc659, n_237, wc660);
  not gc659 (wc660, n_1772);
  and gc658 (wc657, A[2], wc658);
  not gc657 (wc658, n_1304);
  or g2302 (n_246, wc664, wc666, wc667, wc668);
  and gc668 (wc668, n_212, n_241);
  and gc667 (wc667, n_240, n_1812);
  and gc666 (wc666, n_237, n_210);
  and gc665 (wc664, A[3], wc665);
  not gc664 (wc665, n_1304);
  or g2303 (n_2024, B[3], wc669);
  not gc669 (wc669, n_247);
  and g2304 (n_1614, B[4], wc670);
  not gc670 (wc670, n_248);
  or g2305 (n_2025, B[4], wc671);
  not gc671 (wc671, n_248);
  and g2306 (n_2026, B[5], wc672);
  not gc672 (wc672, n_249);
  and g2307 (n_1620, B[6], wc673);
  not gc673 (wc673, n_250);
  or g2308 (n_2027, B[5], wc674);
  not gc674 (wc674, n_249);
  or g2309 (n_2028, B[6], wc675);
  not gc675 (wc675, n_250);
  or g2310 (n_2029, B[1], wc676);
  not gc676 (wc676, n_245);
  and g2311 (n_1608, B[2], wc677);
  not gc677 (wc677, n_246);
  or g2312 (n_2030, B[2], wc678);
  not gc678 (wc678, n_246);
  and g2313 (n_2031, B[1], wc679);
  not gc679 (wc679, n_245);
  and g2314 (n_2032, B[3], wc680);
  not gc680 (wc680, n_247);
  or g2315 (n_2033, B[4], wc681);
  not gc681 (wc681, n_247);
  and g2316 (n_1546, B[5], wc682);
  not gc682 (wc682, n_248);
  or g2317 (n_2034, B[5], wc683);
  not gc683 (wc683, n_248);
  and g2318 (n_1552, B[6], wc684);
  not gc684 (wc684, n_249);
  or g2319 (n_2035, B[6], wc685);
  not gc685 (wc685, n_249);
  or g2320 (n_2036, B[2], wc686);
  not gc686 (wc686, n_245);
  and g2321 (n_1540, B[3], wc687);
  not gc687 (wc687, n_246);
  or g2322 (n_2037, B[3], wc688);
  not gc688 (wc688, n_246);
  and g2323 (n_2038, B[2], wc689);
  not gc689 (wc689, n_245);
  and g2324 (n_2039, B[4], wc690);
  not gc690 (wc690, n_247);
  or g2325 (n_2040, wc691, n_1831);
  not gc691 (wc691, n_251);
  or g2326 (n_2041, wc692, n_43);
  not gc692 (wc692, n_247);
  and g2327 (n_1694, wc693, n_44);
  not gc693 (wc693, n_248);
  or g2328 (n_2042, wc694, n_44);
  not gc694 (wc694, n_248);
  and g2329 (n_2043, wc695, n_45);
  not gc695 (wc695, n_249);
  and g2330 (n_1700, wc696, n_46);
  not gc696 (wc696, n_250);
  or g2331 (n_2044, wc697, n_45);
  not gc697 (wc697, n_249);
  or g2332 (n_2045, wc698, n_46);
  not gc698 (wc698, n_250);
  or g2333 (n_2046, wc699, n_1794);
  not gc699 (wc699, n_245);
  and g2334 (n_1688, wc700, n_42);
  not gc700 (wc700, n_246);
  or g2335 (n_2047, wc701, n_42);
  not gc701 (wc701, n_246);
  and g2336 (n_2048, wc702, n_1794);
  not gc702 (wc702, n_245);
  and g2337 (n_2049, wc703, n_43);
  not gc703 (wc703, n_247);
  and g2338 (n_2050, wc704, n_1831);
  not gc704 (wc704, n_251);
  and g2339 (n_2051, n_2025, wc705);
  not gc705 (wc705, n_1616);
  and g2340 (n_2052, n_2028, wc706);
  not gc706 (wc706, n_1622);
  and g2341 (n_2053, n_2030, wc707);
  not gc707 (wc707, n_1610);
  and g2342 (n_2054, n_2034, wc708);
  not gc708 (wc708, n_1548);
  and g2343 (n_2055, n_2035, wc709);
  not gc709 (wc709, n_250);
  and g2344 (n_2056, n_2037, wc710);
  not gc710 (wc710, n_1542);
  or g2345 (n_2057, n_1552, wc711);
  not gc711 (wc711, n_1562);
  and g2346 (n_2058, n_2042, wc712);
  not gc712 (wc712, n_1696);
  and g2347 (n_2059, n_2045, wc713);
  not gc713 (wc713, n_1702);
  and g2348 (n_2060, n_2047, wc714);
  not gc714 (wc714, n_1690);
  and g2349 (n_2061, wc715, n_1636);
  not gc715 (wc715, n_2051);
  and g2350 (n_2062, wc716, n_1716);
  not gc716 (wc716, n_2058);
  and g2351 (n_2063, wc717, n_2052);
  not gc717 (wc717, n_2061);
  or g2352 (n_2064, n_1649, wc718);
  not gc718 (wc718, n_1641);
  and g2353 (n_2065, n_2055, wc719);
  not gc719 (wc719, n_1565);
  or g2354 (n_2066, n_2057, wc720);
  not gc720 (wc720, n_1567);
  and g2355 (n_2067, wc721, n_2059);
  not gc721 (wc721, n_2062);
  or g2356 (n_2068, n_1729, wc722);
  not gc722 (wc722, n_1721);
  or g2357 (n_2069, n_2050, wc723);
  not gc723 (wc723, n_1734);
  or g2358 (n_2070, n_1653, n_251);
  or g2359 (n_2071, n_1576, n_251);
  and g2360 (n_2072, n_2071, wc724);
  not gc724 (wc724, n_2070);
  or g2361 (QUOTIENT[1], n_286, n_2070);
endmodule

module divide_unsigned_GENERIC(A, B, QUOTIENT);
  input [14:0] A;
  input [6:0] B;
  output [14:0] QUOTIENT;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] QUOTIENT;
  divide_unsigned_GENERIC_REAL g1(.A (A), .B (B), .QUOTIENT (QUOTIENT));
endmodule

module divide_unsigned_267_GENERIC_REAL(A, B, QUOTIENT);
// synthesis_equation "assign QUOTIENT = A / B;"
  input [14:0] A;
  input [6:0] B;
  output [14:0] QUOTIENT;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] QUOTIENT;
  wire n_39, n_40, n_42, n_43, n_44, n_45, n_46, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_56, n_57, n_59;
  wire n_60, n_63, n_64, n_65, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_80;
  wire n_81, n_82, n_85, n_86, n_87, n_88, n_89, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_110, n_111, n_112, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_147, n_150, n_151, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_165, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_192, n_195;
  wire n_196, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_210, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_237, n_240, n_241, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_286, n_302, n_305, n_308, n_310;
  wire n_311, n_312, n_313, n_316, n_317, n_318, n_319, n_322;
  wire n_325, n_327, n_329, n_331, n_332, n_335, n_336, n_342;
  wire n_346, n_348, n_349, n_358, n_360, n_377, n_379, n_381;
  wire n_382, n_383, n_384, n_387, n_388, n_408, n_411, n_413;
  wire n_414, n_415, n_416, n_419, n_420, n_431, n_448, n_450;
  wire n_451, n_452, n_453, n_456, n_457, n_458, n_460, n_468;
  wire n_487, n_489, n_491, n_493, n_494, n_495, n_496, n_498;
  wire n_499, n_500, n_501, n_502, n_505, n_507, n_510, n_512;
  wire n_522, n_535, n_536, n_539, n_541, n_542, n_543, n_544;
  wire n_546, n_547, n_548, n_549, n_550, n_553, n_555, n_558;
  wire n_563, n_570, n_576, n_594, n_596, n_597, n_598, n_599;
  wire n_601, n_602, n_603, n_604, n_605, n_608, n_610, n_613;
  wire n_618, n_625, n_633, n_650, n_652, n_654, n_656, n_657;
  wire n_658, n_659, n_661, n_662, n_663, n_664, n_665, n_667;
  wire n_668, n_671, n_673, n_674, n_675, n_676, n_677, n_679;
  wire n_681, n_684, n_692, n_696, n_698, n_709, n_710, n_713;
  wire n_715, n_716, n_717, n_718, n_720, n_721, n_722, n_723;
  wire n_724, n_726, n_727, n_728, n_729, n_730, n_733, n_735;
  wire n_736, n_739, n_741, n_744, n_747, n_752, n_754, n_759;
  wire n_763, n_765, n_780, n_782, n_783, n_784, n_785, n_787;
  wire n_788, n_789, n_790, n_791, n_793, n_794, n_795, n_796;
  wire n_797, n_800, n_802, n_803, n_806, n_808, n_811, n_814;
  wire n_819, n_821, n_823, n_828, n_832, n_834, n_846, n_848;
  wire n_850, n_852, n_853, n_854, n_855, n_857, n_858, n_859;
  wire n_860, n_861, n_863, n_864, n_865, n_866, n_869, n_871;
  wire n_872, n_875, n_878, n_880, n_883, n_889, n_894, n_898;
  wire n_900, n_914, n_915, n_918, n_920, n_921, n_922, n_923;
  wire n_925, n_926, n_927, n_928, n_929, n_931, n_932, n_933;
  wire n_935, n_937, n_938, n_941, n_943, n_944, n_947, n_949;
  wire n_954, n_957, n_962, n_966, n_971, n_975, n_977, n_998;
  wire n_1000, n_1001, n_1002, n_1003, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1011, n_1012, n_1013, n_1015, n_1017, n_1018, n_1021;
  wire n_1023, n_1024, n_1027, n_1029, n_1034, n_1037, n_1042, n_1047;
  wire n_1054, n_1058, n_1060, n_1075, n_1077, n_1079, n_1081, n_1082;
  wire n_1083, n_1084, n_1086, n_1087, n_1088, n_1089, n_1090, n_1092;
  wire n_1093, n_1094, n_1095, n_1098, n_1100, n_1101, n_1104, n_1107;
  wire n_1109, n_1112, n_1118, n_1123, n_1127, n_1129, n_1143, n_1144;
  wire n_1147, n_1149, n_1150, n_1151, n_1152, n_1154, n_1155, n_1156;
  wire n_1157, n_1158, n_1160, n_1161, n_1162, n_1164, n_1166, n_1167;
  wire n_1170, n_1172, n_1173, n_1176, n_1178, n_1183, n_1186, n_1191;
  wire n_1195, n_1200, n_1204, n_1206, n_1227, n_1229, n_1230, n_1231;
  wire n_1232, n_1234, n_1235, n_1236, n_1237, n_1238, n_1240, n_1241;
  wire n_1242, n_1244, n_1246, n_1247, n_1250, n_1252, n_1253, n_1256;
  wire n_1258, n_1263, n_1266, n_1271, n_1276, n_1283, n_1287, n_1289;
  wire n_1304, n_1306, n_1308, n_1310, n_1311, n_1312, n_1313, n_1315;
  wire n_1316, n_1317, n_1318, n_1319, n_1321, n_1322, n_1323, n_1324;
  wire n_1327, n_1329, n_1330, n_1333, n_1336, n_1338, n_1341, n_1347;
  wire n_1352, n_1356, n_1358, n_1372, n_1373, n_1376, n_1378, n_1379;
  wire n_1380, n_1381, n_1383, n_1384, n_1385, n_1386, n_1387, n_1389;
  wire n_1390, n_1391, n_1393, n_1395, n_1396, n_1399, n_1401, n_1402;
  wire n_1405, n_1407, n_1412, n_1415, n_1420, n_1424, n_1429, n_1433;
  wire n_1435, n_1456, n_1458, n_1459, n_1460, n_1461, n_1463, n_1464;
  wire n_1465, n_1466, n_1467, n_1469, n_1470, n_1471, n_1473, n_1475;
  wire n_1476, n_1479, n_1481, n_1482, n_1485, n_1487, n_1492, n_1495;
  wire n_1500, n_1505, n_1512, n_1516, n_1518, n_1535, n_1540, n_1542;
  wire n_1546, n_1548, n_1552, n_1553, n_1556, n_1558, n_1562, n_1565;
  wire n_1567, n_1576, n_1608, n_1610, n_1614, n_1616, n_1620, n_1622;
  wire n_1625, n_1628, n_1630, n_1634, n_1636, n_1641, n_1649, n_1653;
  wire n_1688, n_1690, n_1694, n_1696, n_1700, n_1702, n_1705, n_1708;
  wire n_1710, n_1714, n_1716, n_1721, n_1729, n_1734, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815;
  wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  wire n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1840;
  wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1865, n_1866;
  wire n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874;
  wire n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882;
  wire n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890;
  wire n_1891, n_1892, n_1893, n_1894, n_1895, n_1898, n_1899, n_1900;
  wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908;
  wire n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916;
  wire n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924;
  wire n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932;
  wire n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1940, n_1941;
  wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
  wire n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957;
  wire n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965;
  wire n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973;
  wire n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1982;
  wire n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990;
  wire n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998;
  wire n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006;
  wire n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014;
  wire n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022;
  wire n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031;
  wire n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039;
  wire n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047;
  wire n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
  wire n_2072;
  not g1 (QUOTIENT[14], n_39);
  nand g11 (QUOTIENT[13], n_56, n_59);
  and g19 (n_82, n_535, n_81);
  and g31 (n_112, n_709, n_111);
  or g46 (QUOTIENT[6], n_151, n_147);
  or g58 (QUOTIENT[4], n_196, n_192);
  or g70 (QUOTIENT[2], n_241, n_237);
  or g82 (QUOTIENT[0], n_286, n_2072);
  xor g84 (n_349, B[0], B[1]);
  nand g2 (n_302, B[0], B[1]);
  nor g87 (n_305, B[1], B[2]);
  nand g88 (n_308, B[1], B[2]);
  nand g90 (n_310, B[2], B[3]);
  nand g92 (n_312, B[3], B[4]);
  nand g13 (n_316, B[4], B[5]);
  nand g15 (n_318, B[5], B[6]);
  nand g95 (n_322, n_308, n_1779);
  nor g96 (n_313, n_310, n_311);
  nor g24 (n_325, n_358, n_311);
  nor g25 (n_319, n_316, n_317);
  nor g99 (n_331, n_360, n_317);
  nand g102 (n_342, n_310, n_1816);
  nand g103 (n_327, n_325, n_322);
  nand g104 (n_332, n_1783, n_327);
  nand g38 (n_336, n_331, B[6]);
  nand g107 (n_346, n_316, n_1829);
  nand g108 (n_335, n_331, n_332);
  nand g109 (n_348, n_329, n_335);
  xnor g50 (n_42, n_322, n_1780);
  xnor g115 (n_43, n_342, n_1782);
  xnor g117 (n_44, n_332, n_1784);
  xnor g120 (n_45, n_346, n_1785);
  nor g126 (n_358, B[2], B[3]);
  nor g36 (n_360, B[4], B[5]);
  nand g158 (n_384, n_379, n_1793);
  nor g159 (n_382, n_381, B[3]);
  nor g160 (n_387, n_383, B[3]);
  nand g165 (n_388, n_387, n_384);
  xnor g175 (n_49, n_377, n_1796);
  xnor g177 (n_51, n_384, n_1832);
  nand g197 (n_416, n_411, n_408);
  nor g198 (n_414, n_413, B[2]);
  nor g199 (n_419, n_415, B[2]);
  nor g200 (n_311, B[3], B[4]);
  nor g201 (n_317, B[5], B[6]);
  nand g205 (n_420, n_419, n_416);
  nand g209 (n_431, n_311, n_317);
  xnor g220 (n_52, n_416, n_1833);
  nand g243 (n_453, n_448, n_1815);
  nor g244 (n_451, n_450, n_42);
  nor g245 (n_456, n_452, n_42);
  nor g246 (n_458, n_43, n_44);
  nor g247 (n_460, n_45, n_46);
  nand g251 (n_457, n_456, n_453);
  nand g255 (n_468, n_458, n_460);
  xnor g266 (n_50, n_377, n_1817);
  xnor g268 (n_53, n_453, n_1834);
  nand g303 (n_502, n_491, n_1798);
  nor g304 (n_496, n_493, n_494);
  nor g307 (n_505, n_498, n_494);
  nor g308 (n_500, n_499, B[5]);
  nor g309 (n_510, n_501, B[5]);
  nand g312 (n_522, n_493, n_1850);
  nand g313 (n_507, n_505, n_502);
  nand g314 (n_512, n_1840, n_507);
  xnor g327 (n_67, n_489, n_1799);
  xnor g329 (n_69, n_502, n_1847);
  xnor g332 (n_72, n_522, n_1851);
  xnor g334 (n_75, n_512, n_1844);
  nand g359 (n_550, n_539, n_536);
  nor g360 (n_544, n_541, n_542);
  nor g363 (n_553, n_546, n_542);
  nor g364 (n_548, n_547, B[4]);
  nor g365 (n_558, n_549, B[4]);
  nand g369 (n_576, n_541, n_1852);
  nand g370 (n_555, n_553, n_550);
  nand g371 (n_563, n_1842, n_555);
  nand g377 (n_570, n_558, n_317);
  xnor g392 (n_70, n_550, n_1848);
  xnor g395 (n_73, n_576, n_1853);
  xnor g397 (n_76, n_563, n_1845);
  nand g423 (n_605, n_594, n_1818);
  nor g424 (n_599, n_596, n_597);
  nor g427 (n_608, n_601, n_597);
  nor g428 (n_603, n_602, n_44);
  nor g429 (n_613, n_604, n_44);
  nand g433 (n_633, n_596, n_1854);
  nand g434 (n_610, n_608, n_605);
  nand g435 (n_618, n_1843, n_610);
  nand g441 (n_625, n_613, n_460);
  xnor g456 (n_68, n_489, n_1819);
  xnor g458 (n_71, n_605, n_1849);
  xnor g461 (n_74, n_633, n_1855);
  xnor g463 (n_77, n_618, n_1846);
  nand g502 (n_668, n_654, n_1801);
  nor g503 (n_659, n_656, n_657);
  nor g506 (n_671, n_661, n_657);
  nor g507 (n_665, n_662, n_663);
  nor g510 (n_679, n_667, n_663);
  nand g513 (n_692, n_656, n_1875);
  nand g514 (n_673, n_671, n_668);
  nand g515 (n_681, n_1865, n_673);
  nor g516 (n_677, n_674, n_675);
  nand g523 (n_696, n_662, n_1893);
  nand g524 (n_684, n_679, n_681);
  nand g525 (n_698, n_675, n_684);
  nand g528 (n_650, n_1889, n_1890);
  xnor g530 (n_91, n_652, n_1802);
  xnor g532 (n_93, n_668, n_1872);
  xnor g535 (n_96, n_692, n_1876);
  xnor g537 (n_99, n_681, n_1881);
  xnor g540 (n_102, n_696, n_1884);
  xnor g542 (n_105, n_698, n_1869);
  nand g569 (n_730, n_713, n_710);
  nor g570 (n_718, n_715, n_716);
  nor g573 (n_733, n_720, n_716);
  nor g574 (n_724, n_721, n_722);
  nor g577 (n_739, n_726, n_722);
  nor g578 (n_728, n_727, B[6]);
  nor g579 (n_741, n_729, B[6]);
  nand g582 (n_759, n_715, n_1877);
  nand g583 (n_735, n_733, n_730);
  nand g584 (n_744, n_1867, n_735);
  nor g592 (n_754, n_1887, n_728);
  nand g593 (n_752, n_739, n_741);
  nand g596 (n_763, n_721, n_1894);
  nand g597 (n_747, n_739, n_744);
  nand g598 (n_765, n_736, n_747);
  nand g604 (n_709, n_754, n_1891);
  xnor g608 (n_94, n_730, n_1873);
  xnor g611 (n_97, n_759, n_1878);
  xnor g613 (n_100, n_744, n_1882);
  xnor g616 (n_103, n_763, n_1885);
  xnor g618 (n_106, n_765, n_1870);
  nand g645 (n_797, n_780, n_1820);
  nor g646 (n_785, n_782, n_783);
  nor g649 (n_800, n_787, n_783);
  nor g650 (n_791, n_788, n_789);
  nor g653 (n_806, n_793, n_789);
  nor g654 (n_795, n_794, n_46);
  nor g655 (n_808, n_796, n_46);
  nand g658 (n_828, n_782, n_1879);
  nand g659 (n_802, n_800, n_797);
  nand g660 (n_811, n_1868, n_802);
  nor g668 (n_821, n_1888, n_795);
  nand g669 (n_819, n_806, n_808);
  nand g672 (n_832, n_788, n_1895);
  nand g673 (n_814, n_806, n_811);
  nand g674 (n_834, n_803, n_814);
  nand g680 (n_823, n_821, n_1892);
  xnor g684 (n_92, n_652, n_1821);
  xnor g686 (n_95, n_797, n_1874);
  xnor g689 (n_98, n_828, n_1880);
  xnor g691 (n_101, n_811, n_1883);
  xnor g694 (n_104, n_832, n_1886);
  xnor g696 (n_107, n_834, n_1871);
  nand g732 (n_866, n_850, n_1804);
  nor g733 (n_855, n_852, n_853);
  nor g736 (n_869, n_857, n_853);
  nor g737 (n_861, n_858, n_859);
  nor g740 (n_875, n_863, n_859);
  nand g744 (n_894, n_852, n_1915);
  nand g745 (n_871, n_869, n_866);
  nand g746 (n_880, n_1903, n_871);
  nor g751 (n_878, n_872, n_865);
  nand g757 (n_898, n_858, n_1935);
  nand g758 (n_883, n_875, n_880);
  nand g759 (n_900, n_872, n_883);
  nand g763 (n_889, n_1929, n_1930);
  xnor g766 (n_123, n_848, n_1805);
  xnor g768 (n_125, n_866, n_1912);
  xnor g771 (n_128, n_894, n_1916);
  xnor g773 (n_131, n_880, n_1921);
  xnor g776 (n_134, n_898, n_1924);
  xnor g778 (n_137, n_900, n_1909);
  nand g812 (n_938, n_918, n_915);
  nor g813 (n_923, n_920, n_921);
  nor g816 (n_941, n_925, n_921);
  nor g817 (n_929, n_926, n_927);
  nor g820 (n_947, n_931, n_927);
  nor g821 (n_935, n_932, n_933);
  nor g824 (n_949, n_937, n_933);
  nand g827 (n_971, n_920, n_1917);
  nand g828 (n_943, n_941, n_938);
  nand g829 (n_954, n_1906, n_943);
  nand g839 (n_962, n_947, n_949);
  nand g842 (n_975, n_926, n_1936);
  nand g843 (n_957, n_947, n_954);
  nand g844 (n_977, n_944, n_957);
  nand g850 (n_966, n_1931, n_1932);
  xnor g855 (n_126, n_938, n_1913);
  xnor g858 (n_129, n_971, n_1918);
  xnor g860 (n_132, n_954, n_1922);
  xnor g863 (n_135, n_975, n_1925);
  xnor g865 (n_138, n_977, n_1910);
  nand g904 (n_1018, n_998, n_1822);
  nor g905 (n_1003, n_1000, n_1001);
  nor g908 (n_1021, n_1005, n_1001);
  nor g909 (n_1009, n_1006, n_1007);
  nor g912 (n_1027, n_1011, n_1007);
  nor g913 (n_1015, n_1012, n_1013);
  nor g916 (n_1029, n_1017, n_1013);
  nand g919 (n_1054, n_1000, n_1919);
  nand g920 (n_1023, n_1021, n_1018);
  nand g921 (n_1034, n_1908, n_1023);
  nand g931 (n_1042, n_1027, n_1029);
  nand g934 (n_1058, n_1006, n_1937);
  nand g935 (n_1037, n_1027, n_1034);
  nand g936 (n_1060, n_1024, n_1037);
  nand g942 (n_1047, n_1933, n_1934);
  nand g945 (n_151, n_1899, n_1938);
  xnor g947 (n_124, n_848, n_1823);
  xnor g949 (n_127, n_1018, n_1914);
  xnor g952 (n_130, n_1054, n_1920);
  xnor g954 (n_133, n_1034, n_1923);
  xnor g957 (n_136, n_1058, n_1926);
  xnor g959 (n_139, n_1060, n_1911);
  nand g1000 (n_1095, n_1079, n_1807);
  nor g1001 (n_1084, n_1081, n_1082);
  nor g1004 (n_1098, n_1086, n_1082);
  nor g1005 (n_1090, n_1087, n_1088);
  nor g1008 (n_1104, n_1092, n_1088);
  nand g1012 (n_1123, n_1081, n_1957);
  nand g1013 (n_1100, n_1098, n_1095);
  nand g1014 (n_1109, n_1945, n_1100);
  nor g1019 (n_1107, n_1101, n_1094);
  nand g1025 (n_1127, n_1087, n_1977);
  nand g1026 (n_1112, n_1104, n_1109);
  nand g1027 (n_1129, n_1101, n_1112);
  nand g1031 (n_1118, n_1971, n_1972);
  xnor g1034 (n_165, n_1077, n_1808);
  xnor g1036 (n_168, n_1095, n_1954);
  xnor g1039 (n_171, n_1123, n_1958);
  xnor g1041 (n_174, n_1109, n_1963);
  xnor g1044 (n_177, n_1127, n_1966);
  xnor g1046 (n_180, n_1129, n_1951);
  nand g1080 (n_1167, n_1147, n_1144);
  nor g1081 (n_1152, n_1149, n_1150);
  nor g1084 (n_1170, n_1154, n_1150);
  nor g1085 (n_1158, n_1155, n_1156);
  nor g1088 (n_1176, n_1160, n_1156);
  nor g1089 (n_1164, n_1161, n_1162);
  nor g1092 (n_1178, n_1166, n_1162);
  nand g1095 (n_1200, n_1149, n_1959);
  nand g1096 (n_1172, n_1170, n_1167);
  nand g1097 (n_1183, n_1948, n_1172);
  nand g1107 (n_1191, n_1176, n_1178);
  nand g1110 (n_1204, n_1155, n_1978);
  nand g1111 (n_1186, n_1176, n_1183);
  nand g1112 (n_1206, n_1173, n_1186);
  nand g1118 (n_1195, n_1973, n_1974);
  xnor g1123 (n_169, n_1167, n_1955);
  xnor g1126 (n_172, n_1200, n_1960);
  xnor g1128 (n_175, n_1183, n_1964);
  xnor g1131 (n_178, n_1204, n_1967);
  xnor g1133 (n_181, n_1206, n_1952);
  nand g1172 (n_1247, n_1227, n_1824);
  nor g1173 (n_1232, n_1229, n_1230);
  nor g1176 (n_1250, n_1234, n_1230);
  nor g1177 (n_1238, n_1235, n_1236);
  nor g1180 (n_1256, n_1240, n_1236);
  nor g1181 (n_1244, n_1241, n_1242);
  nor g1184 (n_1258, n_1246, n_1242);
  nand g1187 (n_1283, n_1229, n_1961);
  nand g1188 (n_1252, n_1250, n_1247);
  nand g1189 (n_1263, n_1950, n_1252);
  nand g1199 (n_1271, n_1256, n_1258);
  nand g1202 (n_1287, n_1235, n_1979);
  nand g1203 (n_1266, n_1256, n_1263);
  nand g1204 (n_1289, n_1253, n_1266);
  nand g1210 (n_1276, n_1975, n_1976);
  nand g1213 (n_196, n_1941, n_1980);
  xnor g1215 (n_167, n_1077, n_1825);
  xnor g1217 (n_170, n_1247, n_1956);
  xnor g1220 (n_173, n_1283, n_1962);
  xnor g1222 (n_176, n_1263, n_1965);
  xnor g1225 (n_179, n_1287, n_1968);
  xnor g1227 (n_182, n_1289, n_1953);
  nand g1268 (n_1324, n_1308, n_1810);
  nor g1269 (n_1313, n_1310, n_1311);
  nor g1272 (n_1327, n_1315, n_1311);
  nor g1273 (n_1319, n_1316, n_1317);
  nor g1276 (n_1333, n_1321, n_1317);
  nand g1280 (n_1352, n_1310, n_1999);
  nand g1281 (n_1329, n_1327, n_1324);
  nand g1282 (n_1338, n_1987, n_1329);
  nor g1287 (n_1336, n_1330, n_1323);
  nand g1293 (n_1356, n_1316, n_2019);
  nand g1294 (n_1341, n_1333, n_1338);
  nand g1295 (n_1358, n_1330, n_1341);
  nand g1299 (n_1347, n_2013, n_2014);
  xnor g1302 (n_210, n_1306, n_1811);
  xnor g1304 (n_213, n_1324, n_1996);
  xnor g1307 (n_216, n_1352, n_2000);
  xnor g1309 (n_219, n_1338, n_2005);
  xnor g1312 (n_222, n_1356, n_2008);
  xnor g1314 (n_225, n_1358, n_1993);
  nand g1348 (n_1396, n_1376, n_1373);
  nor g1349 (n_1381, n_1378, n_1379);
  nor g1352 (n_1399, n_1383, n_1379);
  nor g1353 (n_1387, n_1384, n_1385);
  nor g1356 (n_1405, n_1389, n_1385);
  nor g1357 (n_1393, n_1390, n_1391);
  nor g1360 (n_1407, n_1395, n_1391);
  nand g1363 (n_1429, n_1378, n_2001);
  nand g1364 (n_1401, n_1399, n_1396);
  nand g1365 (n_1412, n_1990, n_1401);
  nand g1375 (n_1420, n_1405, n_1407);
  nand g1378 (n_1433, n_1384, n_2020);
  nand g1379 (n_1415, n_1405, n_1412);
  nand g1380 (n_1435, n_1402, n_1415);
  nand g1386 (n_1424, n_2015, n_2016);
  xnor g1391 (n_214, n_1396, n_1997);
  xnor g1394 (n_217, n_1429, n_2002);
  xnor g1396 (n_220, n_1412, n_2006);
  xnor g1399 (n_223, n_1433, n_2009);
  xnor g1401 (n_226, n_1435, n_1994);
  nand g1440 (n_1476, n_1456, n_1826);
  nor g1441 (n_1461, n_1458, n_1459);
  nor g1444 (n_1479, n_1463, n_1459);
  nor g1445 (n_1467, n_1464, n_1465);
  nor g1448 (n_1485, n_1469, n_1465);
  nor g1449 (n_1473, n_1470, n_1471);
  nor g1452 (n_1487, n_1475, n_1471);
  nand g1455 (n_1512, n_1458, n_2003);
  nand g1456 (n_1481, n_1479, n_1476);
  nand g1457 (n_1492, n_1992, n_1481);
  nand g1467 (n_1500, n_1485, n_1487);
  nand g1470 (n_1516, n_1464, n_2021);
  nand g1471 (n_1495, n_1485, n_1492);
  nand g1472 (n_1518, n_1482, n_1495);
  nand g1478 (n_1505, n_2017, n_2018);
  nand g1481 (n_241, n_1983, n_2022);
  xnor g1483 (n_212, n_1306, n_1827);
  xnor g1485 (n_215, n_1476, n_1998);
  xnor g1488 (n_218, n_1512, n_2004);
  xnor g1490 (n_221, n_1492, n_2007);
  xnor g1493 (n_224, n_1516, n_2010);
  xnor g1495 (n_227, n_1518, n_1995);
  nand g1536 (n_1553, n_1775, n_1813);
  nor g1537 (n_1542, n_2036, n_1540);
  nor g1540 (n_1556, n_2038, n_1540);
  nor g1541 (n_1548, n_2033, n_1546);
  nor g1544 (n_1562, n_2039, n_1546);
  nand g1549 (n_1558, n_1556, n_1553);
  nand g1550 (n_1567, n_2056, n_1558);
  nor g1555 (n_1565, n_2054, n_1552);
  nand g1567 (n_1576, n_2065, n_2066);
  nand g1616 (n_1625, n_1773, n_1774);
  nor g1617 (n_1610, n_2029, n_1608);
  nor g1620 (n_1628, n_2031, n_1608);
  nor g1621 (n_1616, n_2024, n_1614);
  nor g1624 (n_1634, n_2032, n_1614);
  nor g1625 (n_1622, n_2027, n_1620);
  nor g1628 (n_1636, n_2026, n_1620);
  nand g1632 (n_1630, n_1628, n_1625);
  nand g1633 (n_1641, n_2053, n_1630);
  nand g1643 (n_1649, n_1634, n_1636);
  nand g1654 (n_1653, n_2063, n_2064);
  nand g1708 (n_1705, n_1791, n_1828);
  nor g1709 (n_1690, n_2046, n_1688);
  nor g1712 (n_1708, n_2048, n_1688);
  nor g1713 (n_1696, n_2041, n_1694);
  nor g1716 (n_1714, n_2049, n_1694);
  nor g1717 (n_1702, n_2044, n_1700);
  nor g1720 (n_1716, n_2043, n_1700);
  nand g1724 (n_1710, n_1708, n_1705);
  nand g1725 (n_1721, n_2060, n_1710);
  nand g1735 (n_1729, n_1714, n_1716);
  nand g1746 (n_1734, n_2067, n_2068);
  nand g1749 (n_286, n_2040, n_2069);
  or g1781 (n_1758, wc, A[14]);
  not gc (wc, B[0]);
  or g1782 (n_1759, B[6], wc0);
  not gc0 (wc0, n_360);
  xnor g1783 (n_1760, A[14], B[0]);
  or g1784 (n_379, B[1], wc1);
  not gc1 (wc1, A[13]);
  or g1785 (n_377, wc2, A[12]);
  not gc2 (wc2, B[0]);
  and g1786 (n_1761, B[1], wc3);
  not gc3 (wc3, A[13]);
  or g1787 (n_411, B[0], wc4);
  not gc4 (wc4, A[13]);
  and g1788 (n_408, B[0], wc5);
  not gc5 (wc5, A[13]);
  xnor g1789 (n_1762, A[12], B[0]);
  or g1790 (n_491, B[1], wc6);
  not gc6 (wc6, A[11]);
  or g1791 (n_489, wc7, A[10]);
  not gc7 (wc7, B[0]);
  and g1792 (n_1763, B[1], wc8);
  not gc8 (wc8, A[11]);
  or g1793 (n_539, B[0], wc9);
  not gc9 (wc9, A[11]);
  and g1794 (n_536, B[0], wc10);
  not gc10 (wc10, A[11]);
  xnor g1795 (n_1764, A[10], B[0]);
  or g1796 (n_654, B[1], wc11);
  not gc11 (wc11, A[9]);
  or g1797 (n_652, wc12, A[8]);
  not gc12 (wc12, B[0]);
  and g1798 (n_1765, B[1], wc13);
  not gc13 (wc13, A[9]);
  or g1799 (n_713, B[0], wc14);
  not gc14 (wc14, A[9]);
  and g1800 (n_710, B[0], wc15);
  not gc15 (wc15, A[9]);
  xnor g1801 (n_1766, A[8], B[0]);
  or g1802 (n_850, B[1], wc16);
  not gc16 (wc16, A[7]);
  or g1803 (n_848, wc17, A[6]);
  not gc17 (wc17, B[0]);
  and g1804 (n_1767, B[1], wc18);
  not gc18 (wc18, A[7]);
  or g1805 (n_918, B[0], wc19);
  not gc19 (wc19, A[7]);
  and g1806 (n_915, B[0], wc20);
  not gc20 (wc20, A[7]);
  xnor g1807 (n_1768, A[6], B[0]);
  or g1808 (n_1079, B[1], wc21);
  not gc21 (wc21, A[5]);
  or g1809 (n_1077, wc22, A[4]);
  not gc22 (wc22, B[0]);
  and g1810 (n_1769, B[1], wc23);
  not gc23 (wc23, A[5]);
  or g1811 (n_1147, B[0], wc24);
  not gc24 (wc24, A[5]);
  and g1812 (n_1144, B[0], wc25);
  not gc25 (wc25, A[5]);
  xnor g1813 (n_1770, A[4], B[0]);
  or g1814 (n_1308, B[1], wc26);
  not gc26 (wc26, A[3]);
  or g1815 (n_1306, wc27, A[2]);
  not gc27 (wc27, B[0]);
  and g1816 (n_1771, B[1], wc28);
  not gc28 (wc28, A[3]);
  or g1817 (n_1376, B[0], wc29);
  not gc29 (wc29, A[3]);
  and g1818 (n_1373, B[0], wc30);
  not gc30 (wc30, A[3]);
  xnor g1819 (n_1772, A[2], B[0]);
  or g1820 (n_1773, B[0], wc31);
  not gc31 (wc31, A[1]);
  and g1821 (n_1774, B[0], wc32);
  not gc32 (wc32, A[1]);
  or g1822 (n_1775, B[1], wc33);
  not gc33 (wc33, A[1]);
  or g1823 (n_1535, wc34, A[0]);
  not gc34 (wc34, B[0]);
  and g1824 (n_1776, B[1], wc35);
  not gc35 (wc35, A[1]);
  or g1825 (n_1777, B[1], wc36);
  not gc36 (wc36, n_1758);
  or g1826 (n_1778, wc37, n_305);
  not gc37 (wc37, n_308);
  or g1827 (n_1779, n_302, n_305);
  or g1828 (n_1780, n_358, wc38);
  not gc38 (wc38, n_310);
  or g1829 (n_448, wc39, n_349);
  not gc39 (wc39, A[13]);
  and g1830 (n_1781, wc40, n_349);
  not gc40 (wc40, A[13]);
  or g1831 (n_1782, n_311, wc41);
  not gc41 (wc41, n_312);
  and g1832 (n_1783, wc42, n_312);
  not gc42 (wc42, n_313);
  or g1833 (n_1784, n_360, wc43);
  not gc43 (wc43, n_316);
  or g1834 (n_1785, n_317, wc44);
  not gc44 (wc44, n_318);
  and g1835 (n_329, wc45, n_318);
  not gc45 (wc45, n_319);
  or g1836 (n_594, wc46, n_349);
  not gc46 (wc46, A[11]);
  and g1837 (n_1786, wc47, n_349);
  not gc47 (wc47, A[11]);
  or g1838 (n_780, wc48, n_349);
  not gc48 (wc48, A[9]);
  and g1839 (n_1787, wc49, n_349);
  not gc49 (wc49, A[9]);
  or g1840 (n_998, wc50, n_349);
  not gc50 (wc50, A[7]);
  and g1841 (n_1788, wc51, n_349);
  not gc51 (wc51, A[7]);
  or g1842 (n_1227, wc52, n_349);
  not gc52 (wc52, A[5]);
  and g1843 (n_1789, wc53, n_349);
  not gc53 (wc53, A[5]);
  or g1844 (n_1456, wc54, n_349);
  not gc54 (wc54, A[3]);
  and g1845 (n_1790, wc55, n_349);
  not gc55 (wc55, A[3]);
  or g1846 (n_1791, wc56, n_349);
  not gc56 (wc56, A[1]);
  and g1847 (n_1792, wc57, n_349);
  not gc57 (wc57, A[1]);
  or g1848 (n_1793, n_1761, wc58);
  not gc58 (wc58, n_377);
  xor g1849 (n_1794, n_302, n_1778);
  and g1850 (n_1795, B[6], wc59);
  not gc59 (wc59, n_329);
  or g1851 (n_1796, n_1761, wc60);
  not gc60 (wc60, n_379);
  or g1852 (n_1797, n_408, wc61);
  not gc61 (wc61, n_411);
  or g1853 (n_1798, n_1763, wc62);
  not gc62 (wc62, n_489);
  or g1854 (n_1799, n_1763, wc63);
  not gc63 (wc63, n_491);
  or g1855 (n_1800, n_536, wc64);
  not gc64 (wc64, n_539);
  or g1856 (n_1801, n_1765, wc65);
  not gc65 (wc65, n_652);
  or g1857 (n_1802, n_1765, wc66);
  not gc66 (wc66, n_654);
  or g1858 (n_1803, n_710, wc67);
  not gc67 (wc67, n_713);
  or g1859 (n_1804, n_1767, wc68);
  not gc68 (wc68, n_848);
  or g1860 (n_1805, n_1767, wc69);
  not gc69 (wc69, n_850);
  or g1861 (n_1806, n_915, wc70);
  not gc70 (wc70, n_918);
  or g1862 (n_1807, n_1769, wc71);
  not gc71 (wc71, n_1077);
  or g1863 (n_1808, n_1769, wc72);
  not gc72 (wc72, n_1079);
  or g1864 (n_1809, n_1144, wc73);
  not gc73 (wc73, n_1147);
  or g1865 (n_1810, n_1771, wc74);
  not gc74 (wc74, n_1306);
  or g1866 (n_1811, n_1771, wc75);
  not gc75 (wc75, n_1308);
  or g1867 (n_1812, n_1373, wc76);
  not gc76 (wc76, n_1376);
  or g1868 (n_1813, n_1776, wc77);
  not gc77 (wc77, n_1535);
  or g1869 (n_1814, n_1777, wc78);
  not gc78 (wc78, n_358);
  or g1870 (n_1815, n_1781, wc79);
  not gc79 (wc79, n_377);
  or g1871 (n_1816, n_358, wc80);
  not gc80 (wc80, n_322);
  or g1872 (n_1817, n_1781, wc81);
  not gc81 (wc81, n_448);
  or g1873 (n_1818, n_1786, wc82);
  not gc82 (wc82, n_489);
  or g1874 (n_1819, n_1786, wc83);
  not gc83 (wc83, n_594);
  or g1875 (n_1820, n_1787, wc84);
  not gc84 (wc84, n_652);
  or g1876 (n_1821, n_1787, wc85);
  not gc85 (wc85, n_780);
  or g1877 (n_1822, n_1788, wc86);
  not gc86 (wc86, n_848);
  or g1878 (n_1823, n_1788, wc87);
  not gc87 (wc87, n_998);
  or g1879 (n_1824, n_1789, wc88);
  not gc88 (wc88, n_1077);
  or g1880 (n_1825, n_1789, wc89);
  not gc89 (wc89, n_1227);
  or g1881 (n_1826, n_1790, wc90);
  not gc90 (wc90, n_1306);
  or g1882 (n_1827, n_1790, wc91);
  not gc91 (wc91, n_1456);
  or g1883 (n_1828, n_1792, wc92);
  not gc92 (wc92, n_1535);
  or g1884 (n_39, n_1759, n_1814);
  or g1885 (n_1829, n_360, wc93);
  not gc93 (wc93, n_332);
  or g1886 (n_1830, n_336, wc94);
  not gc94 (wc94, n_332);
  or g1887 (n_1831, wc95, n_1795);
  not gc95 (wc95, n_1830);
  or g1888 (n_40, wc96, wc99);
  and gc99 (wc99, A[14], n_39);
  and gc98 (wc96, wc97, wc98);
  not gc97 (wc98, n_1760);
  not gc96 (wc97, n_39);
  xor g1889 (n_46, n_348, B[6]);
  or g1890 (n_381, B[2], wc100);
  not gc100 (wc100, n_40);
  and g1891 (n_383, B[2], wc101);
  not gc101 (wc101, n_40);
  or g1892 (n_413, B[1], wc102);
  not gc102 (wc102, n_40);
  and g1893 (n_415, B[1], wc103);
  not gc103 (wc103, n_40);
  or g1894 (n_450, wc104, n_1794);
  not gc104 (wc104, n_40);
  and g1895 (n_452, wc105, n_1794);
  not gc105 (wc105, n_40);
  or g1896 (n_1832, n_383, wc106);
  not gc106 (wc106, n_381);
  or g1897 (n_1833, n_415, wc107);
  not gc107 (wc107, n_413);
  or g1898 (n_1834, n_452, wc108);
  not gc108 (wc108, n_450);
  or g1899 (n_1835, wc109, n_382);
  not gc109 (wc109, n_388);
  or g1900 (n_1836, wc110, n_414);
  not gc110 (wc110, n_420);
  or g1901 (n_1837, wc111, n_451);
  not gc111 (wc111, n_457);
  or g1902 (n_54, wc112, n_1759);
  not gc112 (wc112, n_1835);
  or g1903 (n_56, wc113, n_431);
  not gc113 (wc113, n_1836);
  or g1904 (n_1838, wc114, n_468);
  not gc114 (wc114, n_1837);
  and g1905 (n_57, n_56, wc115);
  not gc115 (wc115, n_54);
  or g1906 (n_59, n_1831, n_1838);
  and g1907 (n_60, n_59, wc116);
  not gc116 (wc116, n_56);
  or g1908 (QUOTIENT[12], wc117, n_57);
  not gc117 (wc117, n_59);
  or g1909 (n_65, wc118, wc119, wc120, wc121);
  and gc122 (wc121, wc122, n_53);
  not gc121 (wc122, n_59);
  and gc120 (wc120, n_60, n_52);
  and gc119 (wc119, n_57, n_51);
  and gc118 (wc118, n_54, n_40);
  or g1910 (n_63, wc123, wc124, wc126, wc127);
  and gc129 (wc127, wc128, wc129);
  not gc128 (wc129, n_1762);
  not gc127 (wc128, n_59);
  and gc126 (wc126, A[12], n_60);
  and gc125 (wc124, n_57, wc125);
  not gc124 (wc125, n_1762);
  and gc123 (wc123, A[12], n_54);
  or g1911 (n_64, wc130, wc131, wc132, wc133);
  and gc134 (wc133, wc134, n_50);
  not gc133 (wc134, n_59);
  and gc132 (wc132, n_60, n_1797);
  and gc131 (wc131, n_57, n_49);
  and gc130 (wc130, A[13], n_54);
  or g1912 (n_499, B[4], wc135);
  not gc135 (wc135, n_65);
  or g1913 (n_493, B[2], wc136);
  not gc136 (wc136, n_63);
  and g1914 (n_494, B[3], wc137);
  not gc137 (wc137, n_64);
  or g1915 (n_495, B[3], wc138);
  not gc138 (wc138, n_64);
  and g1916 (n_498, B[2], wc139);
  not gc139 (wc139, n_63);
  and g1917 (n_501, B[4], wc140);
  not gc140 (wc140, n_65);
  or g1918 (n_547, B[3], wc141);
  not gc141 (wc141, n_65);
  or g1919 (n_541, B[1], wc142);
  not gc142 (wc142, n_63);
  and g1920 (n_542, B[2], wc143);
  not gc143 (wc143, n_64);
  or g1921 (n_543, B[2], wc144);
  not gc144 (wc144, n_64);
  and g1922 (n_546, B[1], wc145);
  not gc145 (wc145, n_63);
  and g1923 (n_549, B[3], wc146);
  not gc146 (wc146, n_65);
  or g1924 (n_602, wc147, n_43);
  not gc147 (wc147, n_65);
  or g1925 (n_596, wc148, n_1794);
  not gc148 (wc148, n_63);
  and g1926 (n_597, wc149, n_42);
  not gc149 (wc149, n_64);
  or g1927 (n_598, wc150, n_42);
  not gc150 (wc150, n_64);
  and g1928 (n_601, wc151, n_1794);
  not gc151 (wc151, n_63);
  and g1929 (n_604, wc152, n_43);
  not gc152 (wc152, n_65);
  and g1930 (n_1840, n_495, wc153);
  not gc153 (wc153, n_496);
  or g1931 (n_1841, B[6], wc154);
  not gc154 (wc154, n_510);
  and g1932 (n_1842, n_543, wc155);
  not gc155 (wc155, n_544);
  and g1933 (n_1843, n_598, wc156);
  not gc156 (wc156, n_599);
  or g1934 (n_1844, n_501, wc157);
  not gc157 (wc157, n_499);
  or g1935 (n_1845, n_549, wc158);
  not gc158 (wc158, n_547);
  or g1936 (n_1846, n_604, wc159);
  not gc159 (wc159, n_602);
  or g1937 (n_1847, n_498, wc160);
  not gc160 (wc160, n_493);
  or g1938 (n_1848, n_546, wc161);
  not gc161 (wc161, n_541);
  or g1939 (n_1849, n_601, wc162);
  not gc162 (wc162, n_596);
  or g1940 (n_1850, n_498, wc163);
  not gc163 (wc163, n_502);
  or g1941 (n_1851, wc164, n_494);
  not gc164 (wc164, n_495);
  or g1942 (n_1852, n_546, wc165);
  not gc165 (wc165, n_550);
  or g1943 (n_1853, wc166, n_542);
  not gc166 (wc166, n_543);
  or g1944 (n_1854, n_601, wc167);
  not gc167 (wc167, n_605);
  or g1945 (n_1855, wc168, n_597);
  not gc168 (wc168, n_598);
  and g1946 (n_1856, wc169, n_500);
  not gc169 (wc169, B[6]);
  and g1947 (n_1857, n_317, n_548);
  and g1948 (n_1858, n_460, n_603);
  or g1949 (n_1859, n_1841, wc170);
  not gc170 (wc170, n_512);
  or g1950 (n_1860, n_570, wc171);
  not gc171 (wc171, n_563);
  or g1951 (n_1861, n_625, wc172);
  not gc172 (wc172, n_618);
  or g1952 (n_487, wc173, n_1856);
  not gc173 (wc173, n_1859);
  or g1953 (n_535, wc174, n_1857);
  not gc174 (wc174, n_1860);
  or g1954 (n_1862, wc175, n_1858);
  not gc175 (wc175, n_1861);
  or g1955 (n_81, wc176, n_1831);
  not gc176 (wc176, n_1862);
  and g1956 (n_80, wc177, n_487);
  not gc177 (wc177, n_535);
  or g1957 (QUOTIENT[11], wc178, n_535);
  not gc178 (wc178, n_81);
  or g1958 (QUOTIENT[10], n_80, wc179);
  not gc179 (wc179, n_81);
  or g1959 (n_89, wc180, wc182, wc183, wc184);
  and gc185 (wc184, wc185, n_77);
  not gc184 (wc185, n_81);
  and gc183 (wc183, n_76, n_82);
  and gc182 (wc182, n_80, n_75);
  and gc181 (wc180, wc181, n_65);
  not gc180 (wc181, n_487);
  or g1960 (n_87, wc186, wc188, wc189, wc190);
  and gc191 (wc190, wc191, n_71);
  not gc190 (wc191, n_81);
  and gc189 (wc189, n_70, n_82);
  and gc188 (wc188, n_80, n_69);
  and gc187 (wc186, wc187, n_63);
  not gc186 (wc187, n_487);
  or g1961 (n_88, wc192, wc194, wc195, wc196);
  and gc197 (wc196, wc197, n_74);
  not gc196 (wc197, n_81);
  and gc195 (wc195, n_73, n_82);
  and gc194 (wc194, n_80, n_72);
  and gc193 (wc192, wc193, n_64);
  not gc192 (wc193, n_487);
  or g1962 (n_85, wc198, wc200, wc202, wc203);
  and gc205 (wc203, wc204, wc205);
  not gc204 (wc205, n_1764);
  not gc203 (wc204, n_81);
  and gc202 (wc202, A[10], n_82);
  and gc201 (wc200, n_80, wc201);
  not gc200 (wc201, n_1764);
  and gc199 (wc198, A[10], wc199);
  not gc198 (wc199, n_487);
  or g1963 (n_86, wc206, wc208, wc209, wc210);
  and gc211 (wc210, wc211, n_68);
  not gc210 (wc211, n_81);
  and gc209 (wc209, n_1800, n_82);
  and gc208 (wc208, n_80, n_67);
  and gc207 (wc206, A[11], wc207);
  not gc206 (wc207, n_487);
  and g1964 (n_674, B[6], wc212);
  not gc212 (wc212, n_89);
  or g1965 (n_662, B[4], wc213);
  not gc213 (wc213, n_87);
  and g1966 (n_663, B[5], wc214);
  not gc214 (wc214, n_88);
  or g1967 (n_664, B[5], wc215);
  not gc215 (wc215, n_88);
  or g1968 (n_676, B[6], wc216);
  not gc216 (wc216, n_89);
  or g1969 (n_656, B[2], wc217);
  not gc217 (wc217, n_85);
  and g1970 (n_657, B[3], wc218);
  not gc218 (wc218, n_86);
  or g1971 (n_658, B[3], wc219);
  not gc219 (wc219, n_86);
  and g1972 (n_661, B[2], wc220);
  not gc220 (wc220, n_85);
  and g1973 (n_667, B[4], wc221);
  not gc221 (wc221, n_87);
  or g1974 (n_721, B[3], wc222);
  not gc222 (wc222, n_87);
  and g1975 (n_722, B[4], wc223);
  not gc223 (wc223, n_88);
  or g1976 (n_723, B[4], wc224);
  not gc224 (wc224, n_88);
  and g1977 (n_729, B[5], wc225);
  not gc225 (wc225, n_89);
  or g1978 (n_727, B[5], wc226);
  not gc226 (wc226, n_89);
  or g1979 (n_715, B[1], wc227);
  not gc227 (wc227, n_85);
  and g1980 (n_716, B[2], wc228);
  not gc228 (wc228, n_86);
  or g1981 (n_717, B[2], wc229);
  not gc229 (wc229, n_86);
  and g1982 (n_720, B[1], wc230);
  not gc230 (wc230, n_85);
  and g1983 (n_726, B[3], wc231);
  not gc231 (wc231, n_87);
  or g1984 (n_788, wc232, n_43);
  not gc232 (wc232, n_87);
  and g1985 (n_789, wc233, n_44);
  not gc233 (wc233, n_88);
  or g1986 (n_790, wc234, n_44);
  not gc234 (wc234, n_88);
  and g1987 (n_796, wc235, n_45);
  not gc235 (wc235, n_89);
  or g1988 (n_794, wc236, n_45);
  not gc236 (wc236, n_89);
  or g1989 (n_782, wc237, n_1794);
  not gc237 (wc237, n_85);
  and g1990 (n_783, wc238, n_42);
  not gc238 (wc238, n_86);
  or g1991 (n_784, wc239, n_42);
  not gc239 (wc239, n_86);
  and g1992 (n_787, wc240, n_1794);
  not gc240 (wc240, n_85);
  and g1993 (n_793, wc241, n_43);
  not gc241 (wc241, n_87);
  and g1994 (n_675, n_664, wc242);
  not gc242 (wc242, n_665);
  and g1995 (n_1865, n_658, wc243);
  not gc243 (wc243, n_659);
  or g1996 (n_1866, n_674, wc244);
  not gc244 (wc244, n_679);
  and g1997 (n_736, n_723, wc245);
  not gc245 (wc245, n_724);
  and g1998 (n_1867, n_717, wc246);
  not gc246 (wc246, n_718);
  and g1999 (n_803, n_790, wc247);
  not gc247 (wc247, n_791);
  and g2000 (n_1868, n_784, wc248);
  not gc248 (wc248, n_785);
  or g2001 (n_1869, wc249, n_674);
  not gc249 (wc249, n_676);
  or g2002 (n_1870, wc250, n_729);
  not gc250 (wc250, n_727);
  or g2003 (n_1871, wc251, n_796);
  not gc251 (wc251, n_794);
  or g2004 (n_1872, n_661, wc252);
  not gc252 (wc252, n_656);
  or g2005 (n_1873, n_720, wc253);
  not gc253 (wc253, n_715);
  or g2006 (n_1874, n_787, wc254);
  not gc254 (wc254, n_782);
  or g2007 (n_1875, n_661, wc255);
  not gc255 (wc255, n_668);
  or g2008 (n_1876, wc256, n_657);
  not gc256 (wc256, n_658);
  or g2009 (n_1877, n_720, wc257);
  not gc257 (wc257, n_730);
  or g2010 (n_1878, wc258, n_716);
  not gc258 (wc258, n_717);
  or g2011 (n_1879, n_787, wc259);
  not gc259 (wc259, n_797);
  or g2012 (n_1880, wc260, n_783);
  not gc260 (wc260, n_784);
  or g2013 (n_1881, n_667, wc261);
  not gc261 (wc261, n_662);
  or g2014 (n_1882, n_726, wc262);
  not gc262 (wc262, n_721);
  or g2015 (n_1883, n_793, wc263);
  not gc263 (wc263, n_788);
  or g2016 (n_1884, wc264, n_663);
  not gc264 (wc264, n_664);
  or g2017 (n_1885, wc265, n_722);
  not gc265 (wc265, n_723);
  or g2018 (n_1886, wc266, n_789);
  not gc266 (wc266, n_790);
  and g2019 (n_1887, wc267, n_741);
  not gc267 (wc267, n_736);
  and g2020 (n_1888, wc268, n_808);
  not gc268 (wc268, n_803);
  and g2021 (n_1889, n_676, wc269);
  not gc269 (wc269, n_677);
  or g2022 (n_1890, n_1866, wc270);
  not gc270 (wc270, n_681);
  or g2023 (n_1891, n_752, wc271);
  not gc271 (wc271, n_744);
  or g2024 (n_1892, n_819, wc272);
  not gc272 (wc272, n_811);
  or g2025 (n_1893, n_667, wc273);
  not gc273 (wc273, n_681);
  or g2026 (n_1894, n_726, wc274);
  not gc274 (wc274, n_744);
  or g2027 (n_1895, n_793, wc275);
  not gc275 (wc275, n_811);
  or g2028 (n_111, n_1831, wc276);
  not gc276 (wc276, n_823);
  and g2029 (n_110, wc277, n_650);
  not gc277 (wc277, n_709);
  or g2030 (QUOTIENT[9], wc278, n_709);
  not gc278 (wc278, n_111);
  or g2031 (QUOTIENT[8], n_110, wc279);
  not gc279 (wc279, n_111);
  or g2032 (n_121, wc280, wc282, wc283, wc284);
  and gc285 (wc284, wc285, n_107);
  not gc284 (wc285, n_111);
  and gc283 (wc283, n_106, n_112);
  and gc282 (wc282, n_110, n_105);
  and gc281 (wc280, n_89, wc281);
  not gc280 (wc281, n_650);
  or g2033 (n_117, wc286, wc288, wc289, wc290);
  and gc291 (wc290, wc291, n_95);
  not gc290 (wc291, n_111);
  and gc289 (wc289, n_94, n_112);
  and gc288 (wc288, n_110, n_93);
  and gc287 (wc286, n_85, wc287);
  not gc286 (wc287, n_650);
  or g2034 (n_118, wc292, wc294, wc295, wc296);
  and gc297 (wc296, wc297, n_98);
  not gc296 (wc297, n_111);
  and gc295 (wc295, n_97, n_112);
  and gc294 (wc294, n_110, n_96);
  and gc293 (wc292, n_86, wc293);
  not gc292 (wc293, n_650);
  or g2035 (n_119, wc298, wc300, wc301, wc302);
  and gc303 (wc302, wc303, n_101);
  not gc302 (wc303, n_111);
  and gc301 (wc301, n_100, n_112);
  and gc300 (wc300, n_110, n_99);
  and gc299 (wc298, n_87, wc299);
  not gc298 (wc299, n_650);
  or g2036 (n_120, wc304, wc306, wc307, wc308);
  and gc309 (wc308, wc309, n_104);
  not gc308 (wc309, n_111);
  and gc307 (wc307, n_103, n_112);
  and gc306 (wc306, n_110, n_102);
  and gc305 (wc304, n_88, wc305);
  not gc304 (wc305, n_650);
  or g2037 (n_115, wc310, wc312, wc314, wc315);
  and gc317 (wc315, wc316, wc317);
  not gc316 (wc317, n_1766);
  not gc315 (wc316, n_111);
  and gc314 (wc314, A[8], n_112);
  and gc313 (wc312, n_110, wc313);
  not gc312 (wc313, n_1766);
  and gc311 (wc310, A[8], wc311);
  not gc310 (wc311, n_650);
  or g2038 (n_116, wc318, wc320, wc321, wc322);
  and gc323 (wc322, wc323, n_92);
  not gc322 (wc323, n_111);
  and gc321 (wc321, n_1803, n_112);
  and gc320 (wc320, n_110, n_91);
  and gc319 (wc318, A[9], wc319);
  not gc318 (wc319, n_650);
  or g2039 (n_858, B[4], wc324);
  not gc324 (wc324, n_117);
  and g2040 (n_859, B[5], wc325);
  not gc325 (wc325, n_118);
  or g2041 (n_860, B[5], wc326);
  not gc326 (wc326, n_118);
  and g2042 (n_865, B[6], wc327);
  not gc327 (wc327, n_119);
  or g2043 (n_864, B[6], wc328);
  not gc328 (wc328, n_119);
  or g2044 (n_852, B[2], wc329);
  not gc329 (wc329, n_115);
  and g2045 (n_853, B[3], wc330);
  not gc330 (wc330, n_116);
  or g2046 (n_854, B[3], wc331);
  not gc331 (wc331, n_116);
  and g2047 (n_857, B[2], wc332);
  not gc332 (wc332, n_115);
  and g2048 (n_863, B[4], wc333);
  not gc333 (wc333, n_117);
  or g2049 (n_926, B[3], wc334);
  not gc334 (wc334, n_117);
  and g2050 (n_927, B[4], wc335);
  not gc335 (wc335, n_118);
  or g2051 (n_928, B[4], wc336);
  not gc336 (wc336, n_118);
  and g2052 (n_937, B[5], wc337);
  not gc337 (wc337, n_119);
  and g2053 (n_933, B[6], wc338);
  not gc338 (wc338, n_120);
  or g2054 (n_932, B[5], wc339);
  not gc339 (wc339, n_119);
  or g2055 (n_1898, B[6], wc340);
  not gc340 (wc340, n_120);
  or g2056 (n_920, B[1], wc341);
  not gc341 (wc341, n_115);
  and g2057 (n_921, B[2], wc342);
  not gc342 (wc342, n_116);
  or g2058 (n_922, B[2], wc343);
  not gc343 (wc343, n_116);
  and g2059 (n_925, B[1], wc344);
  not gc344 (wc344, n_115);
  and g2060 (n_931, B[3], wc345);
  not gc345 (wc345, n_117);
  or g2061 (n_1899, wc346, n_1831);
  not gc346 (wc346, n_121);
  or g2062 (n_1006, wc347, n_43);
  not gc347 (wc347, n_117);
  and g2063 (n_1007, wc348, n_44);
  not gc348 (wc348, n_118);
  or g2064 (n_1008, wc349, n_44);
  not gc349 (wc349, n_118);
  and g2065 (n_1017, wc350, n_45);
  not gc350 (wc350, n_119);
  and g2066 (n_1013, wc351, n_46);
  not gc351 (wc351, n_120);
  or g2067 (n_1012, wc352, n_45);
  not gc352 (wc352, n_119);
  or g2068 (n_1900, wc353, n_46);
  not gc353 (wc353, n_120);
  or g2069 (n_1000, wc354, n_1794);
  not gc354 (wc354, n_115);
  and g2070 (n_1001, wc355, n_42);
  not gc355 (wc355, n_116);
  or g2071 (n_1002, wc356, n_42);
  not gc356 (wc356, n_116);
  and g2072 (n_1005, wc357, n_1794);
  not gc357 (wc357, n_115);
  and g2073 (n_1011, wc358, n_43);
  not gc358 (wc358, n_117);
  and g2074 (n_1901, wc359, n_1831);
  not gc359 (wc359, n_121);
  and g2075 (n_872, n_860, wc360);
  not gc360 (wc360, n_861);
  and g2076 (n_1902, n_864, wc361);
  not gc361 (wc361, n_120);
  and g2077 (n_1903, n_854, wc362);
  not gc362 (wc362, n_855);
  or g2078 (n_1904, n_865, wc363);
  not gc363 (wc363, n_875);
  and g2079 (n_944, n_928, wc364);
  not gc364 (wc364, n_929);
  and g2080 (n_1905, n_1898, wc365);
  not gc365 (wc365, n_935);
  and g2081 (n_1906, n_922, wc366);
  not gc366 (wc366, n_923);
  and g2082 (n_1024, n_1008, wc367);
  not gc367 (wc367, n_1009);
  and g2083 (n_1907, n_1900, wc368);
  not gc368 (wc368, n_1015);
  and g2084 (n_1908, n_1002, wc369);
  not gc369 (wc369, n_1003);
  or g2085 (n_1909, wc370, n_865);
  not gc370 (wc370, n_864);
  or g2086 (n_1910, wc371, n_937);
  not gc371 (wc371, n_932);
  or g2087 (n_1911, wc372, n_1017);
  not gc372 (wc372, n_1012);
  or g2088 (n_1912, n_857, wc373);
  not gc373 (wc373, n_852);
  or g2089 (n_1913, n_925, wc374);
  not gc374 (wc374, n_920);
  or g2090 (n_1914, n_1005, wc375);
  not gc375 (wc375, n_1000);
  or g2091 (n_1915, n_857, wc376);
  not gc376 (wc376, n_866);
  or g2092 (n_1916, wc377, n_853);
  not gc377 (wc377, n_854);
  or g2093 (n_1917, n_925, wc378);
  not gc378 (wc378, n_938);
  or g2094 (n_1918, wc379, n_921);
  not gc379 (wc379, n_922);
  or g2095 (n_1919, n_1005, wc380);
  not gc380 (wc380, n_1018);
  or g2096 (n_1920, wc381, n_1001);
  not gc381 (wc381, n_1002);
  or g2097 (n_1921, n_863, wc382);
  not gc382 (wc382, n_858);
  or g2098 (n_1922, n_931, wc383);
  not gc383 (wc383, n_926);
  or g2099 (n_1923, n_1011, wc384);
  not gc384 (wc384, n_1006);
  or g2100 (n_1924, wc385, n_859);
  not gc385 (wc385, n_860);
  or g2101 (n_1925, wc386, n_927);
  not gc386 (wc386, n_928);
  or g2102 (n_1926, wc387, n_1007);
  not gc387 (wc387, n_1008);
  and g2103 (n_1927, wc388, n_949);
  not gc388 (wc388, n_944);
  and g2104 (n_1928, wc389, n_1029);
  not gc389 (wc389, n_1024);
  and g2105 (n_1929, n_1902, wc390);
  not gc390 (wc390, n_878);
  or g2106 (n_1930, n_1904, wc391);
  not gc391 (wc391, n_880);
  and g2107 (n_1931, wc392, n_1905);
  not gc392 (wc392, n_1927);
  or g2108 (n_1932, n_962, wc393);
  not gc393 (wc393, n_954);
  and g2109 (n_1933, wc394, n_1907);
  not gc394 (wc394, n_1928);
  or g2110 (n_1934, n_1042, wc395);
  not gc395 (wc395, n_1034);
  or g2111 (n_1935, n_863, wc396);
  not gc396 (wc396, n_880);
  or g2112 (n_1936, n_931, wc397);
  not gc397 (wc397, n_954);
  or g2113 (n_1937, n_1011, wc398);
  not gc398 (wc398, n_1034);
  or g2114 (n_1938, n_1901, wc399);
  not gc399 (wc399, n_1047);
  or g2115 (n_846, n_889, n_121);
  or g2116 (n_914, n_966, n_121);
  and g2117 (n_147, wc400, n_846);
  not gc400 (wc400, n_914);
  and g2118 (n_150, n_914, wc401);
  not gc401 (wc401, n_151);
  or g2119 (QUOTIENT[7], n_151, n_914);
  or g2120 (n_161, wc402, wc404, wc405, wc406);
  and gc406 (wc406, n_139, n_151);
  and gc405 (wc405, n_150, n_138);
  and gc404 (wc404, n_147, n_137);
  and gc403 (wc402, wc403, n_119);
  not gc402 (wc403, n_846);
  or g2121 (n_157, wc407, wc409, wc410, wc411);
  and gc411 (wc411, n_127, n_151);
  and gc410 (wc410, n_150, n_126);
  and gc409 (wc409, n_147, n_125);
  and gc408 (wc407, wc408, n_115);
  not gc407 (wc408, n_846);
  or g2122 (n_158, wc412, wc414, wc415, wc416);
  and gc416 (wc416, n_130, n_151);
  and gc415 (wc415, n_150, n_129);
  and gc414 (wc414, n_147, n_128);
  and gc413 (wc412, wc413, n_116);
  not gc412 (wc413, n_846);
  or g2123 (n_159, wc417, wc419, wc420, wc421);
  and gc421 (wc421, n_133, n_151);
  and gc420 (wc420, n_150, n_132);
  and gc419 (wc419, n_147, n_131);
  and gc418 (wc417, wc418, n_117);
  not gc417 (wc418, n_846);
  or g2124 (n_160, wc422, wc424, wc425, wc426);
  and gc426 (wc426, n_136, n_151);
  and gc425 (wc425, n_150, n_135);
  and gc424 (wc424, n_147, n_134);
  and gc423 (wc422, wc423, n_118);
  not gc422 (wc423, n_846);
  or g2125 (n_155, wc427, wc429, wc431, wc432);
  and gc433 (wc432, wc433, n_151);
  not gc432 (wc433, n_1768);
  and gc431 (wc431, A[6], n_150);
  and gc430 (wc429, n_147, wc430);
  not gc429 (wc430, n_1768);
  and gc428 (wc427, A[6], wc428);
  not gc427 (wc428, n_846);
  or g2126 (n_156, wc434, wc436, wc437, wc438);
  and gc438 (wc438, n_124, n_151);
  and gc437 (wc437, n_150, n_1806);
  and gc436 (wc436, n_147, n_123);
  and gc435 (wc434, A[7], wc435);
  not gc434 (wc435, n_846);
  or g2127 (n_1087, B[4], wc439);
  not gc439 (wc439, n_157);
  and g2128 (n_1088, B[5], wc440);
  not gc440 (wc440, n_158);
  or g2129 (n_1089, B[5], wc441);
  not gc441 (wc441, n_158);
  and g2130 (n_1094, B[6], wc442);
  not gc442 (wc442, n_159);
  or g2131 (n_1093, B[6], wc443);
  not gc443 (wc443, n_159);
  or g2132 (n_1081, B[2], wc444);
  not gc444 (wc444, n_155);
  and g2133 (n_1082, B[3], wc445);
  not gc445 (wc445, n_156);
  or g2134 (n_1083, B[3], wc446);
  not gc446 (wc446, n_156);
  and g2135 (n_1086, B[2], wc447);
  not gc447 (wc447, n_155);
  and g2136 (n_1092, B[4], wc448);
  not gc448 (wc448, n_157);
  or g2137 (n_1155, B[3], wc449);
  not gc449 (wc449, n_157);
  and g2138 (n_1156, B[4], wc450);
  not gc450 (wc450, n_158);
  or g2139 (n_1157, B[4], wc451);
  not gc451 (wc451, n_158);
  and g2140 (n_1166, B[5], wc452);
  not gc452 (wc452, n_159);
  and g2141 (n_1162, B[6], wc453);
  not gc453 (wc453, n_160);
  or g2142 (n_1161, B[5], wc454);
  not gc454 (wc454, n_159);
  or g2143 (n_1940, B[6], wc455);
  not gc455 (wc455, n_160);
  or g2144 (n_1149, B[1], wc456);
  not gc456 (wc456, n_155);
  and g2145 (n_1150, B[2], wc457);
  not gc457 (wc457, n_156);
  or g2146 (n_1151, B[2], wc458);
  not gc458 (wc458, n_156);
  and g2147 (n_1154, B[1], wc459);
  not gc459 (wc459, n_155);
  and g2148 (n_1160, B[3], wc460);
  not gc460 (wc460, n_157);
  or g2149 (n_1941, wc461, n_1831);
  not gc461 (wc461, n_161);
  or g2150 (n_1235, wc462, n_43);
  not gc462 (wc462, n_157);
  and g2151 (n_1236, wc463, n_44);
  not gc463 (wc463, n_158);
  or g2152 (n_1237, wc464, n_44);
  not gc464 (wc464, n_158);
  and g2153 (n_1246, wc465, n_45);
  not gc465 (wc465, n_159);
  and g2154 (n_1242, wc466, n_46);
  not gc466 (wc466, n_160);
  or g2155 (n_1241, wc467, n_45);
  not gc467 (wc467, n_159);
  or g2156 (n_1942, wc468, n_46);
  not gc468 (wc468, n_160);
  or g2157 (n_1229, wc469, n_1794);
  not gc469 (wc469, n_155);
  and g2158 (n_1230, wc470, n_42);
  not gc470 (wc470, n_156);
  or g2159 (n_1231, wc471, n_42);
  not gc471 (wc471, n_156);
  and g2160 (n_1234, wc472, n_1794);
  not gc472 (wc472, n_155);
  and g2161 (n_1240, wc473, n_43);
  not gc473 (wc473, n_157);
  and g2162 (n_1943, wc474, n_1831);
  not gc474 (wc474, n_161);
  and g2163 (n_1101, n_1089, wc475);
  not gc475 (wc475, n_1090);
  and g2164 (n_1944, n_1093, wc476);
  not gc476 (wc476, n_160);
  and g2165 (n_1945, n_1083, wc477);
  not gc477 (wc477, n_1084);
  or g2166 (n_1946, n_1094, wc478);
  not gc478 (wc478, n_1104);
  and g2167 (n_1173, n_1157, wc479);
  not gc479 (wc479, n_1158);
  and g2168 (n_1947, n_1940, wc480);
  not gc480 (wc480, n_1164);
  and g2169 (n_1948, n_1151, wc481);
  not gc481 (wc481, n_1152);
  and g2170 (n_1253, n_1237, wc482);
  not gc482 (wc482, n_1238);
  and g2171 (n_1949, n_1942, wc483);
  not gc483 (wc483, n_1244);
  and g2172 (n_1950, n_1231, wc484);
  not gc484 (wc484, n_1232);
  or g2173 (n_1951, wc485, n_1094);
  not gc485 (wc485, n_1093);
  or g2174 (n_1952, wc486, n_1166);
  not gc486 (wc486, n_1161);
  or g2175 (n_1953, wc487, n_1246);
  not gc487 (wc487, n_1241);
  or g2176 (n_1954, n_1086, wc488);
  not gc488 (wc488, n_1081);
  or g2177 (n_1955, n_1154, wc489);
  not gc489 (wc489, n_1149);
  or g2178 (n_1956, n_1234, wc490);
  not gc490 (wc490, n_1229);
  or g2179 (n_1957, n_1086, wc491);
  not gc491 (wc491, n_1095);
  or g2180 (n_1958, wc492, n_1082);
  not gc492 (wc492, n_1083);
  or g2181 (n_1959, n_1154, wc493);
  not gc493 (wc493, n_1167);
  or g2182 (n_1960, wc494, n_1150);
  not gc494 (wc494, n_1151);
  or g2183 (n_1961, n_1234, wc495);
  not gc495 (wc495, n_1247);
  or g2184 (n_1962, wc496, n_1230);
  not gc496 (wc496, n_1231);
  or g2185 (n_1963, n_1092, wc497);
  not gc497 (wc497, n_1087);
  or g2186 (n_1964, n_1160, wc498);
  not gc498 (wc498, n_1155);
  or g2187 (n_1965, n_1240, wc499);
  not gc499 (wc499, n_1235);
  or g2188 (n_1966, wc500, n_1088);
  not gc500 (wc500, n_1089);
  or g2189 (n_1967, wc501, n_1156);
  not gc501 (wc501, n_1157);
  or g2190 (n_1968, wc502, n_1236);
  not gc502 (wc502, n_1237);
  and g2191 (n_1969, wc503, n_1178);
  not gc503 (wc503, n_1173);
  and g2192 (n_1970, wc504, n_1258);
  not gc504 (wc504, n_1253);
  and g2193 (n_1971, n_1944, wc505);
  not gc505 (wc505, n_1107);
  or g2194 (n_1972, n_1946, wc506);
  not gc506 (wc506, n_1109);
  and g2195 (n_1973, wc507, n_1947);
  not gc507 (wc507, n_1969);
  or g2196 (n_1974, n_1191, wc508);
  not gc508 (wc508, n_1183);
  and g2197 (n_1975, wc509, n_1949);
  not gc509 (wc509, n_1970);
  or g2198 (n_1976, n_1271, wc510);
  not gc510 (wc510, n_1263);
  or g2199 (n_1977, n_1092, wc511);
  not gc511 (wc511, n_1109);
  or g2200 (n_1978, n_1160, wc512);
  not gc512 (wc512, n_1183);
  or g2201 (n_1979, n_1240, wc513);
  not gc513 (wc513, n_1263);
  or g2202 (n_1980, n_1943, wc514);
  not gc514 (wc514, n_1276);
  or g2203 (n_1075, n_1118, n_161);
  or g2204 (n_1143, n_1195, n_161);
  and g2205 (n_192, wc515, n_1075);
  not gc515 (wc515, n_1143);
  and g2206 (n_195, n_1143, wc516);
  not gc516 (wc516, n_196);
  or g2207 (QUOTIENT[5], n_196, n_1143);
  or g2208 (n_206, wc517, wc519, wc520, wc521);
  and gc521 (wc521, n_182, n_196);
  and gc520 (wc520, n_195, n_181);
  and gc519 (wc519, n_192, n_180);
  and gc518 (wc517, wc518, n_159);
  not gc517 (wc518, n_1075);
  or g2209 (n_202, wc522, wc524, wc525, wc526);
  and gc526 (wc526, n_170, n_196);
  and gc525 (wc525, n_195, n_169);
  and gc524 (wc524, n_192, n_168);
  and gc523 (wc522, wc523, n_155);
  not gc522 (wc523, n_1075);
  or g2210 (n_203, wc527, wc529, wc530, wc531);
  and gc531 (wc531, n_173, n_196);
  and gc530 (wc530, n_195, n_172);
  and gc529 (wc529, n_192, n_171);
  and gc528 (wc527, wc528, n_156);
  not gc527 (wc528, n_1075);
  or g2211 (n_204, wc532, wc534, wc535, wc536);
  and gc536 (wc536, n_176, n_196);
  and gc535 (wc535, n_195, n_175);
  and gc534 (wc534, n_192, n_174);
  and gc533 (wc532, wc533, n_157);
  not gc532 (wc533, n_1075);
  or g2212 (n_205, wc537, wc539, wc540, wc541);
  and gc541 (wc541, n_179, n_196);
  and gc540 (wc540, n_195, n_178);
  and gc539 (wc539, n_192, n_177);
  and gc538 (wc537, wc538, n_158);
  not gc537 (wc538, n_1075);
  or g2213 (n_200, wc542, wc544, wc546, wc547);
  and gc548 (wc547, wc548, n_196);
  not gc547 (wc548, n_1770);
  and gc546 (wc546, A[4], n_195);
  and gc545 (wc544, n_192, wc545);
  not gc544 (wc545, n_1770);
  and gc543 (wc542, A[4], wc543);
  not gc542 (wc543, n_1075);
  or g2214 (n_201, wc549, wc551, wc552, wc553);
  and gc553 (wc553, n_167, n_196);
  and gc552 (wc552, n_195, n_1809);
  and gc551 (wc551, n_192, n_165);
  and gc550 (wc549, A[5], wc550);
  not gc549 (wc550, n_1075);
  or g2215 (n_1316, B[4], wc554);
  not gc554 (wc554, n_202);
  and g2216 (n_1317, B[5], wc555);
  not gc555 (wc555, n_203);
  or g2217 (n_1318, B[5], wc556);
  not gc556 (wc556, n_203);
  and g2218 (n_1323, B[6], wc557);
  not gc557 (wc557, n_204);
  or g2219 (n_1322, B[6], wc558);
  not gc558 (wc558, n_204);
  or g2220 (n_1310, B[2], wc559);
  not gc559 (wc559, n_200);
  and g2221 (n_1311, B[3], wc560);
  not gc560 (wc560, n_201);
  or g2222 (n_1312, B[3], wc561);
  not gc561 (wc561, n_201);
  and g2223 (n_1315, B[2], wc562);
  not gc562 (wc562, n_200);
  and g2224 (n_1321, B[4], wc563);
  not gc563 (wc563, n_202);
  or g2225 (n_1384, B[3], wc564);
  not gc564 (wc564, n_202);
  and g2226 (n_1385, B[4], wc565);
  not gc565 (wc565, n_203);
  or g2227 (n_1386, B[4], wc566);
  not gc566 (wc566, n_203);
  and g2228 (n_1395, B[5], wc567);
  not gc567 (wc567, n_204);
  and g2229 (n_1391, B[6], wc568);
  not gc568 (wc568, n_205);
  or g2230 (n_1390, B[5], wc569);
  not gc569 (wc569, n_204);
  or g2231 (n_1982, B[6], wc570);
  not gc570 (wc570, n_205);
  or g2232 (n_1378, B[1], wc571);
  not gc571 (wc571, n_200);
  and g2233 (n_1379, B[2], wc572);
  not gc572 (wc572, n_201);
  or g2234 (n_1380, B[2], wc573);
  not gc573 (wc573, n_201);
  and g2235 (n_1383, B[1], wc574);
  not gc574 (wc574, n_200);
  and g2236 (n_1389, B[3], wc575);
  not gc575 (wc575, n_202);
  or g2237 (n_1983, wc576, n_1831);
  not gc576 (wc576, n_206);
  or g2238 (n_1464, wc577, n_43);
  not gc577 (wc577, n_202);
  and g2239 (n_1465, wc578, n_44);
  not gc578 (wc578, n_203);
  or g2240 (n_1466, wc579, n_44);
  not gc579 (wc579, n_203);
  and g2241 (n_1475, wc580, n_45);
  not gc580 (wc580, n_204);
  and g2242 (n_1471, wc581, n_46);
  not gc581 (wc581, n_205);
  or g2243 (n_1470, wc582, n_45);
  not gc582 (wc582, n_204);
  or g2244 (n_1984, wc583, n_46);
  not gc583 (wc583, n_205);
  or g2245 (n_1458, wc584, n_1794);
  not gc584 (wc584, n_200);
  and g2246 (n_1459, wc585, n_42);
  not gc585 (wc585, n_201);
  or g2247 (n_1460, wc586, n_42);
  not gc586 (wc586, n_201);
  and g2248 (n_1463, wc587, n_1794);
  not gc587 (wc587, n_200);
  and g2249 (n_1469, wc588, n_43);
  not gc588 (wc588, n_202);
  and g2250 (n_1985, wc589, n_1831);
  not gc589 (wc589, n_206);
  and g2251 (n_1330, n_1318, wc590);
  not gc590 (wc590, n_1319);
  and g2252 (n_1986, n_1322, wc591);
  not gc591 (wc591, n_205);
  and g2253 (n_1987, n_1312, wc592);
  not gc592 (wc592, n_1313);
  or g2254 (n_1988, n_1323, wc593);
  not gc593 (wc593, n_1333);
  and g2255 (n_1402, n_1386, wc594);
  not gc594 (wc594, n_1387);
  and g2256 (n_1989, n_1982, wc595);
  not gc595 (wc595, n_1393);
  and g2257 (n_1990, n_1380, wc596);
  not gc596 (wc596, n_1381);
  and g2258 (n_1482, n_1466, wc597);
  not gc597 (wc597, n_1467);
  and g2259 (n_1991, n_1984, wc598);
  not gc598 (wc598, n_1473);
  and g2260 (n_1992, n_1460, wc599);
  not gc599 (wc599, n_1461);
  or g2261 (n_1993, wc600, n_1323);
  not gc600 (wc600, n_1322);
  or g2262 (n_1994, wc601, n_1395);
  not gc601 (wc601, n_1390);
  or g2263 (n_1995, wc602, n_1475);
  not gc602 (wc602, n_1470);
  or g2264 (n_1996, n_1315, wc603);
  not gc603 (wc603, n_1310);
  or g2265 (n_1997, n_1383, wc604);
  not gc604 (wc604, n_1378);
  or g2266 (n_1998, n_1463, wc605);
  not gc605 (wc605, n_1458);
  or g2267 (n_1999, n_1315, wc606);
  not gc606 (wc606, n_1324);
  or g2268 (n_2000, wc607, n_1311);
  not gc607 (wc607, n_1312);
  or g2269 (n_2001, n_1383, wc608);
  not gc608 (wc608, n_1396);
  or g2270 (n_2002, wc609, n_1379);
  not gc609 (wc609, n_1380);
  or g2271 (n_2003, n_1463, wc610);
  not gc610 (wc610, n_1476);
  or g2272 (n_2004, wc611, n_1459);
  not gc611 (wc611, n_1460);
  or g2273 (n_2005, n_1321, wc612);
  not gc612 (wc612, n_1316);
  or g2274 (n_2006, n_1389, wc613);
  not gc613 (wc613, n_1384);
  or g2275 (n_2007, n_1469, wc614);
  not gc614 (wc614, n_1464);
  or g2276 (n_2008, wc615, n_1317);
  not gc615 (wc615, n_1318);
  or g2277 (n_2009, wc616, n_1385);
  not gc616 (wc616, n_1386);
  or g2278 (n_2010, wc617, n_1465);
  not gc617 (wc617, n_1466);
  and g2279 (n_2011, wc618, n_1407);
  not gc618 (wc618, n_1402);
  and g2280 (n_2012, wc619, n_1487);
  not gc619 (wc619, n_1482);
  and g2281 (n_2013, n_1986, wc620);
  not gc620 (wc620, n_1336);
  or g2282 (n_2014, n_1988, wc621);
  not gc621 (wc621, n_1338);
  and g2283 (n_2015, wc622, n_1989);
  not gc622 (wc622, n_2011);
  or g2284 (n_2016, n_1420, wc623);
  not gc623 (wc623, n_1412);
  and g2285 (n_2017, wc624, n_1991);
  not gc624 (wc624, n_2012);
  or g2286 (n_2018, n_1500, wc625);
  not gc625 (wc625, n_1492);
  or g2287 (n_2019, n_1321, wc626);
  not gc626 (wc626, n_1338);
  or g2288 (n_2020, n_1389, wc627);
  not gc627 (wc627, n_1412);
  or g2289 (n_2021, n_1469, wc628);
  not gc628 (wc628, n_1492);
  or g2290 (n_2022, n_1985, wc629);
  not gc629 (wc629, n_1505);
  or g2291 (n_1304, n_1347, n_206);
  or g2292 (n_1372, n_1424, n_206);
  and g2293 (n_237, wc630, n_1304);
  not gc630 (wc630, n_1372);
  and g2294 (n_240, n_1372, wc631);
  not gc631 (wc631, n_241);
  or g2295 (QUOTIENT[3], n_241, n_1372);
  or g2296 (n_251, wc632, wc634, wc635, wc636);
  and gc636 (wc636, n_227, n_241);
  and gc635 (wc635, n_240, n_226);
  and gc634 (wc634, n_237, n_225);
  and gc633 (wc632, wc633, n_204);
  not gc632 (wc633, n_1304);
  or g2297 (n_247, wc637, wc639, wc640, wc641);
  and gc641 (wc641, n_215, n_241);
  and gc640 (wc640, n_240, n_214);
  and gc639 (wc639, n_237, n_213);
  and gc638 (wc637, wc638, n_200);
  not gc637 (wc638, n_1304);
  or g2298 (n_248, wc642, wc644, wc645, wc646);
  and gc646 (wc646, n_218, n_241);
  and gc645 (wc645, n_240, n_217);
  and gc644 (wc644, n_237, n_216);
  and gc643 (wc642, wc643, n_201);
  not gc642 (wc643, n_1304);
  or g2299 (n_249, wc647, wc649, wc650, wc651);
  and gc651 (wc651, n_221, n_241);
  and gc650 (wc650, n_240, n_220);
  and gc649 (wc649, n_237, n_219);
  and gc648 (wc647, wc648, n_202);
  not gc647 (wc648, n_1304);
  or g2300 (n_250, wc652, wc654, wc655, wc656);
  and gc656 (wc656, n_224, n_241);
  and gc655 (wc655, n_240, n_223);
  and gc654 (wc654, n_237, n_222);
  and gc653 (wc652, wc653, n_203);
  not gc652 (wc653, n_1304);
  or g2301 (n_245, wc657, wc659, wc661, wc662);
  and gc663 (wc662, wc663, n_241);
  not gc662 (wc663, n_1772);
  and gc661 (wc661, A[2], n_240);
  and gc660 (wc659, n_237, wc660);
  not gc659 (wc660, n_1772);
  and gc658 (wc657, A[2], wc658);
  not gc657 (wc658, n_1304);
  or g2302 (n_246, wc664, wc666, wc667, wc668);
  and gc668 (wc668, n_212, n_241);
  and gc667 (wc667, n_240, n_1812);
  and gc666 (wc666, n_237, n_210);
  and gc665 (wc664, A[3], wc665);
  not gc664 (wc665, n_1304);
  or g2303 (n_2024, B[3], wc669);
  not gc669 (wc669, n_247);
  and g2304 (n_1614, B[4], wc670);
  not gc670 (wc670, n_248);
  or g2305 (n_2025, B[4], wc671);
  not gc671 (wc671, n_248);
  and g2306 (n_2026, B[5], wc672);
  not gc672 (wc672, n_249);
  and g2307 (n_1620, B[6], wc673);
  not gc673 (wc673, n_250);
  or g2308 (n_2027, B[5], wc674);
  not gc674 (wc674, n_249);
  or g2309 (n_2028, B[6], wc675);
  not gc675 (wc675, n_250);
  or g2310 (n_2029, B[1], wc676);
  not gc676 (wc676, n_245);
  and g2311 (n_1608, B[2], wc677);
  not gc677 (wc677, n_246);
  or g2312 (n_2030, B[2], wc678);
  not gc678 (wc678, n_246);
  and g2313 (n_2031, B[1], wc679);
  not gc679 (wc679, n_245);
  and g2314 (n_2032, B[3], wc680);
  not gc680 (wc680, n_247);
  or g2315 (n_2033, B[4], wc681);
  not gc681 (wc681, n_247);
  and g2316 (n_1546, B[5], wc682);
  not gc682 (wc682, n_248);
  or g2317 (n_2034, B[5], wc683);
  not gc683 (wc683, n_248);
  and g2318 (n_1552, B[6], wc684);
  not gc684 (wc684, n_249);
  or g2319 (n_2035, B[6], wc685);
  not gc685 (wc685, n_249);
  or g2320 (n_2036, B[2], wc686);
  not gc686 (wc686, n_245);
  and g2321 (n_1540, B[3], wc687);
  not gc687 (wc687, n_246);
  or g2322 (n_2037, B[3], wc688);
  not gc688 (wc688, n_246);
  and g2323 (n_2038, B[2], wc689);
  not gc689 (wc689, n_245);
  and g2324 (n_2039, B[4], wc690);
  not gc690 (wc690, n_247);
  or g2325 (n_2040, wc691, n_1831);
  not gc691 (wc691, n_251);
  or g2326 (n_2041, wc692, n_43);
  not gc692 (wc692, n_247);
  and g2327 (n_1694, wc693, n_44);
  not gc693 (wc693, n_248);
  or g2328 (n_2042, wc694, n_44);
  not gc694 (wc694, n_248);
  and g2329 (n_2043, wc695, n_45);
  not gc695 (wc695, n_249);
  and g2330 (n_1700, wc696, n_46);
  not gc696 (wc696, n_250);
  or g2331 (n_2044, wc697, n_45);
  not gc697 (wc697, n_249);
  or g2332 (n_2045, wc698, n_46);
  not gc698 (wc698, n_250);
  or g2333 (n_2046, wc699, n_1794);
  not gc699 (wc699, n_245);
  and g2334 (n_1688, wc700, n_42);
  not gc700 (wc700, n_246);
  or g2335 (n_2047, wc701, n_42);
  not gc701 (wc701, n_246);
  and g2336 (n_2048, wc702, n_1794);
  not gc702 (wc702, n_245);
  and g2337 (n_2049, wc703, n_43);
  not gc703 (wc703, n_247);
  and g2338 (n_2050, wc704, n_1831);
  not gc704 (wc704, n_251);
  and g2339 (n_2051, n_2025, wc705);
  not gc705 (wc705, n_1616);
  and g2340 (n_2052, n_2028, wc706);
  not gc706 (wc706, n_1622);
  and g2341 (n_2053, n_2030, wc707);
  not gc707 (wc707, n_1610);
  and g2342 (n_2054, n_2034, wc708);
  not gc708 (wc708, n_1548);
  and g2343 (n_2055, n_2035, wc709);
  not gc709 (wc709, n_250);
  and g2344 (n_2056, n_2037, wc710);
  not gc710 (wc710, n_1542);
  or g2345 (n_2057, n_1552, wc711);
  not gc711 (wc711, n_1562);
  and g2346 (n_2058, n_2042, wc712);
  not gc712 (wc712, n_1696);
  and g2347 (n_2059, n_2045, wc713);
  not gc713 (wc713, n_1702);
  and g2348 (n_2060, n_2047, wc714);
  not gc714 (wc714, n_1690);
  and g2349 (n_2061, wc715, n_1636);
  not gc715 (wc715, n_2051);
  and g2350 (n_2062, wc716, n_1716);
  not gc716 (wc716, n_2058);
  and g2351 (n_2063, wc717, n_2052);
  not gc717 (wc717, n_2061);
  or g2352 (n_2064, n_1649, wc718);
  not gc718 (wc718, n_1641);
  and g2353 (n_2065, n_2055, wc719);
  not gc719 (wc719, n_1565);
  or g2354 (n_2066, n_2057, wc720);
  not gc720 (wc720, n_1567);
  and g2355 (n_2067, wc721, n_2059);
  not gc721 (wc721, n_2062);
  or g2356 (n_2068, n_1729, wc722);
  not gc722 (wc722, n_1721);
  or g2357 (n_2069, n_2050, wc723);
  not gc723 (wc723, n_1734);
  or g2358 (n_2070, n_1653, n_251);
  or g2359 (n_2071, n_1576, n_251);
  and g2360 (n_2072, n_2071, wc724);
  not gc724 (wc724, n_2070);
  or g2361 (QUOTIENT[1], n_286, n_2070);
endmodule

module divide_unsigned_267_GENERIC(A, B, QUOTIENT);
  input [14:0] A;
  input [6:0] B;
  output [14:0] QUOTIENT;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] QUOTIENT;
  divide_unsigned_267_GENERIC_REAL g1(.A (A), .B (B), .QUOTIENT
       (QUOTIENT));
endmodule

module remainder_unsigned_GENERIC_REAL(A, B, REMAINDER);
// synthesis_equation "assign REMAINDER = A % B;"
  input [14:0] A;
  input [6:0] B;
  output [14:0] REMAINDER;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] REMAINDER;
  wire n_32, n_34, n_36, n_37, n_38, n_39, n_40, n_43;
  wire n_44, n_45, n_46, n_47, n_48, n_50, n_51, n_53;
  wire n_54, n_56, n_57, n_58, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_73;
  wire n_74, n_75, n_77, n_78, n_79, n_80, n_81, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_102, n_104, n_105, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_120, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_147, n_150, n_151, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_165, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_192, n_195;
  wire n_196, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_210, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_237, n_240, n_241, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_255, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_282, n_285, n_286, n_295;
  wire n_298, n_301, n_303, n_304, n_305, n_306, n_309, n_310;
  wire n_311, n_312, n_315, n_318, n_320, n_322, n_324, n_325;
  wire n_328, n_329, n_335, n_339, n_341, n_342, n_351, n_353;
  wire n_370, n_372, n_374, n_375, n_376, n_377, n_380, n_381;
  wire n_401, n_404, n_406, n_407, n_408, n_409, n_412, n_413;
  wire n_424, n_441, n_443, n_444, n_445, n_446, n_449, n_450;
  wire n_451, n_453, n_461, n_480, n_482, n_484, n_486, n_487;
  wire n_488, n_489, n_491, n_492, n_493, n_494, n_495, n_498;
  wire n_500, n_503, n_505, n_515, n_528, n_529, n_532, n_534;
  wire n_535, n_536, n_537, n_539, n_540, n_541, n_542, n_543;
  wire n_546, n_548, n_551, n_556, n_563, n_569, n_587, n_589;
  wire n_590, n_591, n_592, n_594, n_595, n_596, n_597, n_598;
  wire n_601, n_603, n_606, n_611, n_618, n_626, n_643, n_645;
  wire n_647, n_649, n_650, n_651, n_652, n_654, n_655, n_656;
  wire n_657, n_658, n_660, n_661, n_664, n_666, n_667, n_668;
  wire n_669, n_670, n_672, n_674, n_677, n_685, n_689, n_691;
  wire n_702, n_703, n_706, n_708, n_709, n_710, n_711, n_713;
  wire n_714, n_715, n_716, n_717, n_719, n_720, n_721, n_722;
  wire n_723, n_726, n_728, n_729, n_732, n_734, n_737, n_740;
  wire n_745, n_747, n_752, n_756, n_758, n_773, n_775, n_776;
  wire n_777, n_778, n_780, n_781, n_782, n_783, n_784, n_786;
  wire n_787, n_788, n_789, n_790, n_793, n_795, n_796, n_799;
  wire n_801, n_804, n_807, n_812, n_814, n_816, n_821, n_825;
  wire n_827, n_839, n_841, n_843, n_845, n_846, n_847, n_848;
  wire n_850, n_851, n_852, n_853, n_854, n_856, n_857, n_858;
  wire n_859, n_862, n_864, n_865, n_868, n_871, n_873, n_876;
  wire n_882, n_887, n_891, n_893, n_907, n_908, n_911, n_913;
  wire n_914, n_915, n_916, n_918, n_919, n_920, n_921, n_922;
  wire n_924, n_925, n_926, n_928, n_930, n_931, n_934, n_936;
  wire n_937, n_940, n_942, n_947, n_950, n_955, n_959, n_964;
  wire n_968, n_970, n_991, n_993, n_994, n_995, n_996, n_998;
  wire n_999, n_1000, n_1001, n_1002, n_1004, n_1005, n_1006, n_1008;
  wire n_1010, n_1011, n_1014, n_1016, n_1017, n_1020, n_1022, n_1027;
  wire n_1030, n_1035, n_1040, n_1047, n_1051, n_1053, n_1068, n_1070;
  wire n_1072, n_1074, n_1075, n_1076, n_1077, n_1079, n_1080, n_1081;
  wire n_1082, n_1083, n_1085, n_1086, n_1087, n_1088, n_1091, n_1093;
  wire n_1094, n_1097, n_1100, n_1102, n_1105, n_1111, n_1116, n_1120;
  wire n_1122, n_1136, n_1137, n_1140, n_1142, n_1143, n_1144, n_1145;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1153, n_1154, n_1155;
  wire n_1157, n_1159, n_1160, n_1163, n_1165, n_1166, n_1169, n_1171;
  wire n_1176, n_1179, n_1184, n_1188, n_1193, n_1197, n_1199, n_1220;
  wire n_1222, n_1223, n_1224, n_1225, n_1227, n_1228, n_1229, n_1230;
  wire n_1231, n_1233, n_1234, n_1235, n_1237, n_1239, n_1240, n_1243;
  wire n_1245, n_1246, n_1249, n_1251, n_1256, n_1259, n_1264, n_1269;
  wire n_1276, n_1280, n_1282, n_1297, n_1299, n_1301, n_1303, n_1304;
  wire n_1305, n_1306, n_1308, n_1309, n_1310, n_1311, n_1312, n_1314;
  wire n_1315, n_1316, n_1317, n_1320, n_1322, n_1323, n_1326, n_1329;
  wire n_1331, n_1334, n_1340, n_1345, n_1349, n_1351, n_1365, n_1366;
  wire n_1369, n_1371, n_1372, n_1373, n_1374, n_1376, n_1377, n_1378;
  wire n_1379, n_1380, n_1382, n_1383, n_1384, n_1386, n_1388, n_1389;
  wire n_1392, n_1394, n_1395, n_1398, n_1400, n_1405, n_1408, n_1413;
  wire n_1417, n_1422, n_1426, n_1428, n_1449, n_1451, n_1452, n_1453;
  wire n_1454, n_1456, n_1457, n_1458, n_1459, n_1460, n_1462, n_1463;
  wire n_1464, n_1466, n_1468, n_1469, n_1472, n_1474, n_1475, n_1478;
  wire n_1480, n_1485, n_1488, n_1493, n_1498, n_1505, n_1509, n_1511;
  wire n_1526, n_1528, n_1530, n_1532, n_1533, n_1534, n_1535, n_1537;
  wire n_1538, n_1539, n_1540, n_1541, n_1543, n_1544, n_1545, n_1546;
  wire n_1549, n_1551, n_1552, n_1555, n_1558, n_1560, n_1563, n_1569;
  wire n_1574, n_1578, n_1580, n_1594, n_1595, n_1598, n_1600, n_1601;
  wire n_1602, n_1603, n_1605, n_1606, n_1607, n_1608, n_1609, n_1611;
  wire n_1612, n_1613, n_1615, n_1617, n_1618, n_1621, n_1623, n_1624;
  wire n_1627, n_1629, n_1634, n_1637, n_1642, n_1646, n_1651, n_1655;
  wire n_1657, n_1678, n_1680, n_1681, n_1682, n_1683, n_1685, n_1686;
  wire n_1687, n_1688, n_1689, n_1691, n_1692, n_1693, n_1695, n_1697;
  wire n_1698, n_1701, n_1703, n_1704, n_1707, n_1709, n_1714, n_1717;
  wire n_1722, n_1727, n_1734, n_1738, n_1740, n_1750, n_1751, n_1752;
  wire n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760;
  wire n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768;
  wire n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832;
  wire n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840;
  wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864;
  wire n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872;
  wire n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880;
  wire n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888;
  wire n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896;
  wire n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904;
  wire n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912;
  wire n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920;
  wire n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928;
  wire n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936;
  wire n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960;
  wire n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976;
  wire n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984;
  wire n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992;
  wire n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000;
  wire n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016;
  wire n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024;
  wire n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032;
  wire n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040;
  wire n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048;
  assign REMAINDER[7] = 1'b0;
  assign REMAINDER[8] = 1'b0;
  assign REMAINDER[9] = 1'b0;
  assign REMAINDER[10] = 1'b0;
  assign REMAINDER[11] = 1'b0;
  assign REMAINDER[12] = 1'b0;
  assign REMAINDER[13] = 1'b0;
  assign REMAINDER[14] = 1'b0;
  and g19 (n_75, n_528, n_74);
  and g31 (n_105, n_702, n_104);
  xor g84 (n_342, B[0], B[1]);
  nand g2 (n_295, B[0], B[1]);
  nor g87 (n_298, B[1], B[2]);
  nand g88 (n_301, B[1], B[2]);
  nand g90 (n_303, B[2], B[3]);
  nand g92 (n_305, B[3], B[4]);
  nand g13 (n_309, B[4], B[5]);
  nand g15 (n_311, B[5], B[6]);
  nand g95 (n_315, n_301, n_1769);
  nor g96 (n_306, n_303, n_304);
  nor g24 (n_318, n_351, n_304);
  nor g25 (n_312, n_309, n_310);
  nor g99 (n_324, n_353, n_310);
  nand g102 (n_335, n_303, n_1807);
  nand g103 (n_320, n_318, n_315);
  nand g104 (n_325, n_1773, n_320);
  nand g38 (n_329, n_324, B[6]);
  nand g107 (n_339, n_309, n_1821);
  nand g108 (n_328, n_324, n_325);
  nand g109 (n_341, n_322, n_328);
  xnor g50 (n_36, n_315, n_1770);
  xnor g115 (n_37, n_335, n_1772);
  xnor g117 (n_38, n_325, n_1774);
  xnor g120 (n_39, n_339, n_1775);
  nor g126 (n_351, B[2], B[3]);
  nor g36 (n_353, B[4], B[5]);
  nand g158 (n_377, n_372, n_1782);
  nor g159 (n_375, n_374, B[3]);
  nor g160 (n_380, n_376, B[3]);
  nand g165 (n_381, n_380, n_377);
  xnor g175 (n_43, n_370, n_1785);
  xnor g177 (n_45, n_377, n_1824);
  nand g197 (n_409, n_404, n_401);
  nor g198 (n_407, n_406, B[2]);
  nor g199 (n_412, n_408, B[2]);
  nor g200 (n_304, B[3], B[4]);
  nor g201 (n_310, B[5], B[6]);
  nand g205 (n_413, n_412, n_409);
  nand g209 (n_424, n_304, n_310);
  xnor g220 (n_46, n_409, n_1825);
  nand g243 (n_446, n_441, n_1806);
  nor g244 (n_444, n_443, n_36);
  nor g245 (n_449, n_445, n_36);
  nor g246 (n_451, n_37, n_38);
  nor g247 (n_453, n_39, n_40);
  nand g251 (n_450, n_449, n_446);
  nand g255 (n_461, n_451, n_453);
  xnor g266 (n_44, n_370, n_1808);
  xnor g268 (n_47, n_446, n_1826);
  nand g303 (n_495, n_484, n_1787);
  nor g304 (n_489, n_486, n_487);
  nor g307 (n_498, n_491, n_487);
  nor g308 (n_493, n_492, B[5]);
  nor g309 (n_503, n_494, B[5]);
  nand g312 (n_515, n_486, n_1841);
  nand g313 (n_500, n_498, n_495);
  nand g314 (n_505, n_1831, n_500);
  xnor g327 (n_60, n_482, n_1788);
  xnor g329 (n_62, n_495, n_1838);
  xnor g332 (n_65, n_515, n_1842);
  xnor g334 (n_68, n_505, n_1835);
  nand g359 (n_543, n_532, n_529);
  nor g360 (n_537, n_534, n_535);
  nor g363 (n_546, n_539, n_535);
  nor g364 (n_541, n_540, B[4]);
  nor g365 (n_551, n_542, B[4]);
  nand g369 (n_569, n_534, n_1843);
  nand g370 (n_548, n_546, n_543);
  nand g371 (n_556, n_1833, n_548);
  nand g377 (n_563, n_551, n_310);
  xnor g392 (n_63, n_543, n_1839);
  xnor g395 (n_66, n_569, n_1844);
  xnor g397 (n_69, n_556, n_1836);
  nand g423 (n_598, n_587, n_1809);
  nor g424 (n_592, n_589, n_590);
  nor g427 (n_601, n_594, n_590);
  nor g428 (n_596, n_595, n_38);
  nor g429 (n_606, n_597, n_38);
  nand g433 (n_626, n_589, n_1845);
  nand g434 (n_603, n_601, n_598);
  nand g435 (n_611, n_1834, n_603);
  nand g441 (n_618, n_606, n_453);
  xnor g456 (n_61, n_482, n_1810);
  xnor g458 (n_64, n_598, n_1840);
  xnor g461 (n_67, n_626, n_1846);
  xnor g463 (n_70, n_611, n_1837);
  nand g502 (n_661, n_647, n_1790);
  nor g503 (n_652, n_649, n_650);
  nor g506 (n_664, n_654, n_650);
  nor g507 (n_658, n_655, n_656);
  nor g510 (n_672, n_660, n_656);
  nand g513 (n_685, n_649, n_1864);
  nand g514 (n_666, n_664, n_661);
  nand g515 (n_674, n_1854, n_666);
  nor g516 (n_670, n_667, n_668);
  nand g523 (n_689, n_655, n_1882);
  nand g524 (n_677, n_672, n_674);
  nand g525 (n_691, n_668, n_677);
  nand g528 (n_643, n_1878, n_1879);
  xnor g530 (n_83, n_645, n_1791);
  xnor g532 (n_85, n_661, n_1861);
  xnor g535 (n_88, n_685, n_1865);
  xnor g537 (n_91, n_674, n_1870);
  xnor g540 (n_94, n_689, n_1873);
  xnor g542 (n_97, n_691, n_1858);
  nand g569 (n_723, n_706, n_703);
  nor g570 (n_711, n_708, n_709);
  nor g573 (n_726, n_713, n_709);
  nor g574 (n_717, n_714, n_715);
  nor g577 (n_732, n_719, n_715);
  nor g578 (n_721, n_720, B[6]);
  nor g579 (n_734, n_722, B[6]);
  nand g582 (n_752, n_708, n_1866);
  nand g583 (n_728, n_726, n_723);
  nand g584 (n_737, n_1856, n_728);
  nor g592 (n_747, n_1876, n_721);
  nand g593 (n_745, n_732, n_734);
  nand g596 (n_756, n_714, n_1883);
  nand g597 (n_740, n_732, n_737);
  nand g598 (n_758, n_729, n_740);
  nand g604 (n_702, n_747, n_1880);
  xnor g608 (n_86, n_723, n_1862);
  xnor g611 (n_89, n_752, n_1867);
  xnor g613 (n_92, n_737, n_1871);
  xnor g616 (n_95, n_756, n_1874);
  xnor g618 (n_98, n_758, n_1859);
  nand g645 (n_790, n_773, n_1811);
  nor g646 (n_778, n_775, n_776);
  nor g649 (n_793, n_780, n_776);
  nor g650 (n_784, n_781, n_782);
  nor g653 (n_799, n_786, n_782);
  nor g654 (n_788, n_787, n_40);
  nor g655 (n_801, n_789, n_40);
  nand g658 (n_821, n_775, n_1868);
  nand g659 (n_795, n_793, n_790);
  nand g660 (n_804, n_1857, n_795);
  nor g668 (n_814, n_1877, n_788);
  nand g669 (n_812, n_799, n_801);
  nand g672 (n_825, n_781, n_1884);
  nand g673 (n_807, n_799, n_804);
  nand g674 (n_827, n_796, n_807);
  nand g680 (n_816, n_814, n_1881);
  xnor g684 (n_84, n_645, n_1812);
  xnor g686 (n_87, n_790, n_1863);
  xnor g689 (n_90, n_821, n_1869);
  xnor g691 (n_93, n_804, n_1872);
  xnor g694 (n_96, n_825, n_1875);
  xnor g696 (n_99, n_827, n_1860);
  nand g732 (n_859, n_843, n_1793);
  nor g733 (n_848, n_845, n_846);
  nor g736 (n_862, n_850, n_846);
  nor g737 (n_854, n_851, n_852);
  nor g740 (n_868, n_856, n_852);
  nand g744 (n_887, n_845, n_1902);
  nand g745 (n_864, n_862, n_859);
  nand g746 (n_873, n_1890, n_864);
  nor g751 (n_871, n_865, n_858);
  nand g757 (n_891, n_851, n_1922);
  nand g758 (n_876, n_868, n_873);
  nand g759 (n_893, n_865, n_876);
  nand g763 (n_882, n_1916, n_1917);
  xnor g766 (n_120, n_841, n_1794);
  xnor g768 (n_123, n_859, n_1899);
  xnor g771 (n_126, n_887, n_1903);
  xnor g773 (n_129, n_873, n_1908);
  xnor g776 (n_132, n_891, n_1911);
  xnor g778 (n_135, n_893, n_1896);
  nand g812 (n_931, n_911, n_908);
  nor g813 (n_916, n_913, n_914);
  nor g816 (n_934, n_918, n_914);
  nor g817 (n_922, n_919, n_920);
  nor g820 (n_940, n_924, n_920);
  nor g821 (n_928, n_925, n_926);
  nor g824 (n_942, n_930, n_926);
  nand g827 (n_964, n_913, n_1904);
  nand g828 (n_936, n_934, n_931);
  nand g829 (n_947, n_1893, n_936);
  nand g839 (n_955, n_940, n_942);
  nand g842 (n_968, n_919, n_1923);
  nand g843 (n_950, n_940, n_947);
  nand g844 (n_970, n_937, n_950);
  nand g850 (n_959, n_1918, n_1919);
  xnor g855 (n_124, n_931, n_1900);
  xnor g858 (n_127, n_964, n_1905);
  xnor g860 (n_130, n_947, n_1909);
  xnor g863 (n_133, n_968, n_1912);
  xnor g865 (n_136, n_970, n_1897);
  nand g904 (n_1011, n_991, n_1813);
  nor g905 (n_996, n_993, n_994);
  nor g908 (n_1014, n_998, n_994);
  nor g909 (n_1002, n_999, n_1000);
  nor g912 (n_1020, n_1004, n_1000);
  nor g913 (n_1008, n_1005, n_1006);
  nor g916 (n_1022, n_1010, n_1006);
  nand g919 (n_1047, n_993, n_1906);
  nand g920 (n_1016, n_1014, n_1011);
  nand g921 (n_1027, n_1895, n_1016);
  nand g931 (n_1035, n_1020, n_1022);
  nand g934 (n_1051, n_999, n_1924);
  nand g935 (n_1030, n_1020, n_1027);
  nand g936 (n_1053, n_1017, n_1030);
  nand g942 (n_1040, n_1920, n_1921);
  nand g945 (n_151, n_1886, n_1925);
  xnor g947 (n_122, n_841, n_1814);
  xnor g949 (n_125, n_1011, n_1901);
  xnor g952 (n_128, n_1047, n_1907);
  xnor g954 (n_131, n_1027, n_1910);
  xnor g957 (n_134, n_1051, n_1913);
  xnor g959 (n_137, n_1053, n_1898);
  nand g1000 (n_1088, n_1072, n_1796);
  nor g1001 (n_1077, n_1074, n_1075);
  nor g1004 (n_1091, n_1079, n_1075);
  nor g1005 (n_1083, n_1080, n_1081);
  nor g1008 (n_1097, n_1085, n_1081);
  nand g1012 (n_1116, n_1074, n_1943);
  nand g1013 (n_1093, n_1091, n_1088);
  nand g1014 (n_1102, n_1931, n_1093);
  nor g1019 (n_1100, n_1094, n_1087);
  nand g1025 (n_1120, n_1080, n_1963);
  nand g1026 (n_1105, n_1097, n_1102);
  nand g1027 (n_1122, n_1094, n_1105);
  nand g1031 (n_1111, n_1957, n_1958);
  xnor g1034 (n_165, n_1070, n_1797);
  xnor g1036 (n_168, n_1088, n_1940);
  xnor g1039 (n_171, n_1116, n_1944);
  xnor g1041 (n_174, n_1102, n_1949);
  xnor g1044 (n_177, n_1120, n_1952);
  xnor g1046 (n_180, n_1122, n_1937);
  nand g1080 (n_1160, n_1140, n_1137);
  nor g1081 (n_1145, n_1142, n_1143);
  nor g1084 (n_1163, n_1147, n_1143);
  nor g1085 (n_1151, n_1148, n_1149);
  nor g1088 (n_1169, n_1153, n_1149);
  nor g1089 (n_1157, n_1154, n_1155);
  nor g1092 (n_1171, n_1159, n_1155);
  nand g1095 (n_1193, n_1142, n_1945);
  nand g1096 (n_1165, n_1163, n_1160);
  nand g1097 (n_1176, n_1934, n_1165);
  nand g1107 (n_1184, n_1169, n_1171);
  nand g1110 (n_1197, n_1148, n_1964);
  nand g1111 (n_1179, n_1169, n_1176);
  nand g1112 (n_1199, n_1166, n_1179);
  nand g1118 (n_1188, n_1959, n_1960);
  xnor g1123 (n_169, n_1160, n_1941);
  xnor g1126 (n_172, n_1193, n_1946);
  xnor g1128 (n_175, n_1176, n_1950);
  xnor g1131 (n_178, n_1197, n_1953);
  xnor g1133 (n_181, n_1199, n_1938);
  nand g1172 (n_1240, n_1220, n_1815);
  nor g1173 (n_1225, n_1222, n_1223);
  nor g1176 (n_1243, n_1227, n_1223);
  nor g1177 (n_1231, n_1228, n_1229);
  nor g1180 (n_1249, n_1233, n_1229);
  nor g1181 (n_1237, n_1234, n_1235);
  nor g1184 (n_1251, n_1239, n_1235);
  nand g1187 (n_1276, n_1222, n_1947);
  nand g1188 (n_1245, n_1243, n_1240);
  nand g1189 (n_1256, n_1936, n_1245);
  nand g1199 (n_1264, n_1249, n_1251);
  nand g1202 (n_1280, n_1228, n_1965);
  nand g1203 (n_1259, n_1249, n_1256);
  nand g1204 (n_1282, n_1246, n_1259);
  nand g1210 (n_1269, n_1961, n_1962);
  nand g1213 (n_196, n_1927, n_1966);
  xnor g1215 (n_167, n_1070, n_1816);
  xnor g1217 (n_170, n_1240, n_1942);
  xnor g1220 (n_173, n_1276, n_1948);
  xnor g1222 (n_176, n_1256, n_1951);
  xnor g1225 (n_179, n_1280, n_1954);
  xnor g1227 (n_182, n_1282, n_1939);
  nand g1268 (n_1317, n_1301, n_1799);
  nor g1269 (n_1306, n_1303, n_1304);
  nor g1272 (n_1320, n_1308, n_1304);
  nor g1273 (n_1312, n_1309, n_1310);
  nor g1276 (n_1326, n_1314, n_1310);
  nand g1280 (n_1345, n_1303, n_1984);
  nand g1281 (n_1322, n_1320, n_1317);
  nand g1282 (n_1331, n_1972, n_1322);
  nor g1287 (n_1329, n_1323, n_1316);
  nand g1293 (n_1349, n_1309, n_2004);
  nand g1294 (n_1334, n_1326, n_1331);
  nand g1295 (n_1351, n_1323, n_1334);
  nand g1299 (n_1340, n_1998, n_1999);
  xnor g1302 (n_210, n_1299, n_1800);
  xnor g1304 (n_213, n_1317, n_1981);
  xnor g1307 (n_216, n_1345, n_1985);
  xnor g1309 (n_219, n_1331, n_1990);
  xnor g1312 (n_222, n_1349, n_1993);
  xnor g1314 (n_225, n_1351, n_1978);
  nand g1348 (n_1389, n_1369, n_1366);
  nor g1349 (n_1374, n_1371, n_1372);
  nor g1352 (n_1392, n_1376, n_1372);
  nor g1353 (n_1380, n_1377, n_1378);
  nor g1356 (n_1398, n_1382, n_1378);
  nor g1357 (n_1386, n_1383, n_1384);
  nor g1360 (n_1400, n_1388, n_1384);
  nand g1363 (n_1422, n_1371, n_1986);
  nand g1364 (n_1394, n_1392, n_1389);
  nand g1365 (n_1405, n_1975, n_1394);
  nand g1375 (n_1413, n_1398, n_1400);
  nand g1378 (n_1426, n_1377, n_2005);
  nand g1379 (n_1408, n_1398, n_1405);
  nand g1380 (n_1428, n_1395, n_1408);
  nand g1386 (n_1417, n_2000, n_2001);
  xnor g1391 (n_214, n_1389, n_1982);
  xnor g1394 (n_217, n_1422, n_1987);
  xnor g1396 (n_220, n_1405, n_1991);
  xnor g1399 (n_223, n_1426, n_1994);
  xnor g1401 (n_226, n_1428, n_1979);
  nand g1440 (n_1469, n_1449, n_1817);
  nor g1441 (n_1454, n_1451, n_1452);
  nor g1444 (n_1472, n_1456, n_1452);
  nor g1445 (n_1460, n_1457, n_1458);
  nor g1448 (n_1478, n_1462, n_1458);
  nor g1449 (n_1466, n_1463, n_1464);
  nor g1452 (n_1480, n_1468, n_1464);
  nand g1455 (n_1505, n_1451, n_1988);
  nand g1456 (n_1474, n_1472, n_1469);
  nand g1457 (n_1485, n_1977, n_1474);
  nand g1467 (n_1493, n_1478, n_1480);
  nand g1470 (n_1509, n_1457, n_2006);
  nand g1471 (n_1488, n_1478, n_1485);
  nand g1472 (n_1511, n_1475, n_1488);
  nand g1478 (n_1498, n_2002, n_2003);
  nand g1481 (n_241, n_1968, n_2007);
  xnor g1483 (n_212, n_1299, n_1818);
  xnor g1485 (n_215, n_1469, n_1983);
  xnor g1488 (n_218, n_1505, n_1989);
  xnor g1490 (n_221, n_1485, n_1992);
  xnor g1493 (n_224, n_1509, n_1995);
  xnor g1495 (n_227, n_1511, n_1980);
  nand g1536 (n_1546, n_1530, n_1802);
  nor g1537 (n_1535, n_1532, n_1533);
  nor g1540 (n_1549, n_1537, n_1533);
  nor g1541 (n_1541, n_1538, n_1539);
  nor g1544 (n_1555, n_1543, n_1539);
  nand g1548 (n_1574, n_1532, n_2019);
  nand g1549 (n_1551, n_1549, n_1546);
  nand g1550 (n_1560, n_2013, n_1551);
  nor g1555 (n_1558, n_1552, n_1545);
  nand g1561 (n_1578, n_1538, n_2045);
  nand g1562 (n_1563, n_1555, n_1560);
  nand g1563 (n_1580, n_1552, n_1563);
  nand g1567 (n_1569, n_2039, n_2040);
  xnor g1570 (n_255, n_1528, n_1803);
  xnor g1572 (n_258, n_1546, n_2020);
  xnor g1575 (n_261, n_1574, n_2021);
  xnor g1577 (n_264, n_1560, n_2022);
  xnor g1580 (n_267, n_1578, n_2023);
  xnor g1582 (n_270, n_1580, n_2024);
  nand g1616 (n_1618, n_1598, n_1595);
  nor g1617 (n_1603, n_1600, n_1601);
  nor g1620 (n_1621, n_1605, n_1601);
  nor g1621 (n_1609, n_1606, n_1607);
  nor g1624 (n_1627, n_1611, n_1607);
  nor g1625 (n_1615, n_1612, n_1613);
  nor g1628 (n_1629, n_1617, n_1613);
  nand g1631 (n_1651, n_1600, n_2025);
  nand g1632 (n_1623, n_1621, n_1618);
  nand g1633 (n_1634, n_2016, n_1623);
  nand g1643 (n_1642, n_1627, n_1629);
  nand g1646 (n_1655, n_1606, n_2046);
  nand g1647 (n_1637, n_1627, n_1634);
  nand g1648 (n_1657, n_1624, n_1637);
  nand g1654 (n_1646, n_2041, n_2042);
  xnor g1659 (n_259, n_1618, n_2026);
  xnor g1662 (n_262, n_1651, n_2027);
  xnor g1664 (n_265, n_1634, n_2028);
  xnor g1667 (n_268, n_1655, n_2029);
  xnor g1669 (n_271, n_1657, n_2030);
  nand g1708 (n_1698, n_1678, n_1819);
  nor g1709 (n_1683, n_1680, n_1681);
  nor g1712 (n_1701, n_1685, n_1681);
  nor g1713 (n_1689, n_1686, n_1687);
  nor g1716 (n_1707, n_1691, n_1687);
  nor g1717 (n_1695, n_1692, n_1693);
  nor g1720 (n_1709, n_1697, n_1693);
  nand g1723 (n_1734, n_1680, n_2031);
  nand g1724 (n_1703, n_1701, n_1698);
  nand g1725 (n_1714, n_2018, n_1703);
  nand g1735 (n_1722, n_1707, n_1709);
  nand g1738 (n_1738, n_1686, n_2047);
  nand g1739 (n_1717, n_1707, n_1714);
  nand g1740 (n_1740, n_1704, n_1717);
  nand g1746 (n_1727, n_2043, n_2044);
  nand g1749 (n_286, n_2009, n_2048);
  xnor g1751 (n_257, n_1528, n_1820);
  xnor g1753 (n_260, n_1698, n_2032);
  xnor g1756 (n_263, n_1734, n_2033);
  xnor g1758 (n_266, n_1714, n_2034);
  xnor g1761 (n_269, n_1738, n_2035);
  xnor g1763 (n_272, n_1740, n_2036);
  or g1781 (n_1750, wc, A[14]);
  not gc (wc, B[0]);
  or g1782 (n_1751, B[6], wc0);
  not gc0 (wc0, n_353);
  xnor g1783 (n_1752, A[14], B[0]);
  or g1784 (n_372, B[1], wc1);
  not gc1 (wc1, A[13]);
  or g1785 (n_370, wc2, A[12]);
  not gc2 (wc2, B[0]);
  and g1786 (n_1753, B[1], wc3);
  not gc3 (wc3, A[13]);
  or g1787 (n_404, B[0], wc4);
  not gc4 (wc4, A[13]);
  and g1788 (n_401, B[0], wc5);
  not gc5 (wc5, A[13]);
  xnor g1789 (n_1754, A[12], B[0]);
  or g1790 (n_484, B[1], wc6);
  not gc6 (wc6, A[11]);
  or g1791 (n_482, wc7, A[10]);
  not gc7 (wc7, B[0]);
  and g1792 (n_1755, B[1], wc8);
  not gc8 (wc8, A[11]);
  or g1793 (n_532, B[0], wc9);
  not gc9 (wc9, A[11]);
  and g1794 (n_529, B[0], wc10);
  not gc10 (wc10, A[11]);
  xnor g1795 (n_1756, A[10], B[0]);
  or g1796 (n_647, B[1], wc11);
  not gc11 (wc11, A[9]);
  or g1797 (n_645, wc12, A[8]);
  not gc12 (wc12, B[0]);
  and g1798 (n_1757, B[1], wc13);
  not gc13 (wc13, A[9]);
  or g1799 (n_706, B[0], wc14);
  not gc14 (wc14, A[9]);
  and g1800 (n_703, B[0], wc15);
  not gc15 (wc15, A[9]);
  xnor g1801 (n_1758, A[8], B[0]);
  or g1802 (n_843, B[1], wc16);
  not gc16 (wc16, A[7]);
  or g1803 (n_841, wc17, A[6]);
  not gc17 (wc17, B[0]);
  and g1804 (n_1759, B[1], wc18);
  not gc18 (wc18, A[7]);
  or g1805 (n_911, B[0], wc19);
  not gc19 (wc19, A[7]);
  and g1806 (n_908, B[0], wc20);
  not gc20 (wc20, A[7]);
  xnor g1807 (n_1760, A[6], B[0]);
  or g1808 (n_1072, B[1], wc21);
  not gc21 (wc21, A[5]);
  or g1809 (n_1070, wc22, A[4]);
  not gc22 (wc22, B[0]);
  and g1810 (n_1761, B[1], wc23);
  not gc23 (wc23, A[5]);
  or g1811 (n_1140, B[0], wc24);
  not gc24 (wc24, A[5]);
  and g1812 (n_1137, B[0], wc25);
  not gc25 (wc25, A[5]);
  xnor g1813 (n_1762, A[4], B[0]);
  or g1814 (n_1301, B[1], wc26);
  not gc26 (wc26, A[3]);
  or g1815 (n_1299, wc27, A[2]);
  not gc27 (wc27, B[0]);
  and g1816 (n_1763, B[1], wc28);
  not gc28 (wc28, A[3]);
  or g1817 (n_1369, B[0], wc29);
  not gc29 (wc29, A[3]);
  and g1818 (n_1366, B[0], wc30);
  not gc30 (wc30, A[3]);
  xnor g1819 (n_1764, A[2], B[0]);
  or g1820 (n_1530, B[1], wc31);
  not gc31 (wc31, A[1]);
  or g1821 (n_1528, wc32, A[0]);
  not gc32 (wc32, B[0]);
  and g1822 (n_1765, B[1], wc33);
  not gc33 (wc33, A[1]);
  or g1823 (n_1598, B[0], wc34);
  not gc34 (wc34, A[1]);
  and g1824 (n_1595, B[0], wc35);
  not gc35 (wc35, A[1]);
  xnor g1825 (n_1766, A[0], B[0]);
  or g1826 (n_1767, B[1], wc36);
  not gc36 (wc36, n_1750);
  or g1827 (n_1768, wc37, n_298);
  not gc37 (wc37, n_301);
  or g1828 (n_1769, n_295, n_298);
  or g1829 (n_1770, n_351, wc38);
  not gc38 (wc38, n_303);
  or g1830 (n_441, wc39, n_342);
  not gc39 (wc39, A[13]);
  and g1831 (n_1771, wc40, n_342);
  not gc40 (wc40, A[13]);
  or g1832 (n_1772, n_304, wc41);
  not gc41 (wc41, n_305);
  and g1833 (n_1773, wc42, n_305);
  not gc42 (wc42, n_306);
  or g1834 (n_1774, n_353, wc43);
  not gc43 (wc43, n_309);
  or g1835 (n_1775, n_310, wc44);
  not gc44 (wc44, n_311);
  and g1836 (n_322, wc45, n_311);
  not gc45 (wc45, n_312);
  or g1837 (n_587, wc46, n_342);
  not gc46 (wc46, A[11]);
  and g1838 (n_1776, wc47, n_342);
  not gc47 (wc47, A[11]);
  or g1839 (n_773, wc48, n_342);
  not gc48 (wc48, A[9]);
  and g1840 (n_1777, wc49, n_342);
  not gc49 (wc49, A[9]);
  or g1841 (n_991, wc50, n_342);
  not gc50 (wc50, A[7]);
  and g1842 (n_1778, wc51, n_342);
  not gc51 (wc51, A[7]);
  or g1843 (n_1220, wc52, n_342);
  not gc52 (wc52, A[5]);
  and g1844 (n_1779, wc53, n_342);
  not gc53 (wc53, A[5]);
  or g1845 (n_1449, wc54, n_342);
  not gc54 (wc54, A[3]);
  and g1846 (n_1780, wc55, n_342);
  not gc55 (wc55, A[3]);
  or g1847 (n_1678, wc56, n_342);
  not gc56 (wc56, A[1]);
  and g1848 (n_1781, wc57, n_342);
  not gc57 (wc57, A[1]);
  or g1849 (n_1782, n_1753, wc58);
  not gc58 (wc58, n_370);
  xor g1850 (n_1783, n_295, n_1768);
  and g1851 (n_1784, B[6], wc59);
  not gc59 (wc59, n_322);
  or g1852 (n_1785, n_1753, wc60);
  not gc60 (wc60, n_372);
  or g1853 (n_1786, n_401, wc61);
  not gc61 (wc61, n_404);
  or g1854 (n_1787, n_1755, wc62);
  not gc62 (wc62, n_482);
  or g1855 (n_1788, n_1755, wc63);
  not gc63 (wc63, n_484);
  or g1856 (n_1789, n_529, wc64);
  not gc64 (wc64, n_532);
  or g1857 (n_1790, n_1757, wc65);
  not gc65 (wc65, n_645);
  or g1858 (n_1791, n_1757, wc66);
  not gc66 (wc66, n_647);
  or g1859 (n_1792, n_703, wc67);
  not gc67 (wc67, n_706);
  or g1860 (n_1793, n_1759, wc68);
  not gc68 (wc68, n_841);
  or g1861 (n_1794, n_1759, wc69);
  not gc69 (wc69, n_843);
  or g1862 (n_1795, n_908, wc70);
  not gc70 (wc70, n_911);
  or g1863 (n_1796, n_1761, wc71);
  not gc71 (wc71, n_1070);
  or g1864 (n_1797, n_1761, wc72);
  not gc72 (wc72, n_1072);
  or g1865 (n_1798, n_1137, wc73);
  not gc73 (wc73, n_1140);
  or g1866 (n_1799, n_1763, wc74);
  not gc74 (wc74, n_1299);
  or g1867 (n_1800, n_1763, wc75);
  not gc75 (wc75, n_1301);
  or g1868 (n_1801, n_1366, wc76);
  not gc76 (wc76, n_1369);
  or g1869 (n_1802, n_1765, wc77);
  not gc77 (wc77, n_1528);
  or g1870 (n_1803, n_1765, wc78);
  not gc78 (wc78, n_1530);
  or g1871 (n_1804, n_1595, wc79);
  not gc79 (wc79, n_1598);
  or g1872 (n_1805, n_1767, wc80);
  not gc80 (wc80, n_351);
  or g1873 (n_1806, n_1771, wc81);
  not gc81 (wc81, n_370);
  or g1874 (n_1807, n_351, wc82);
  not gc82 (wc82, n_315);
  or g1875 (n_1808, n_1771, wc83);
  not gc83 (wc83, n_441);
  or g1876 (n_1809, n_1776, wc84);
  not gc84 (wc84, n_482);
  or g1877 (n_1810, n_1776, wc85);
  not gc85 (wc85, n_587);
  or g1878 (n_1811, n_1777, wc86);
  not gc86 (wc86, n_645);
  or g1879 (n_1812, n_1777, wc87);
  not gc87 (wc87, n_773);
  or g1880 (n_1813, n_1778, wc88);
  not gc88 (wc88, n_841);
  or g1881 (n_1814, n_1778, wc89);
  not gc89 (wc89, n_991);
  or g1882 (n_1815, n_1779, wc90);
  not gc90 (wc90, n_1070);
  or g1883 (n_1816, n_1779, wc91);
  not gc91 (wc91, n_1220);
  or g1884 (n_1817, n_1780, wc92);
  not gc92 (wc92, n_1299);
  or g1885 (n_1818, n_1780, wc93);
  not gc93 (wc93, n_1449);
  or g1886 (n_1819, n_1781, wc94);
  not gc94 (wc94, n_1528);
  or g1887 (n_1820, n_1781, wc95);
  not gc95 (wc95, n_1678);
  or g1888 (n_32, n_1751, n_1805);
  or g1889 (n_1821, n_353, wc96);
  not gc96 (wc96, n_325);
  or g1890 (n_1822, n_329, wc97);
  not gc97 (wc97, n_325);
  or g1891 (n_1823, wc98, n_1784);
  not gc98 (wc98, n_1822);
  or g1892 (n_34, wc99, wc102);
  and gc102 (wc102, A[14], n_32);
  and gc101 (wc99, wc100, wc101);
  not gc100 (wc101, n_1752);
  not gc99 (wc100, n_32);
  xor g1893 (n_40, n_341, B[6]);
  or g1894 (n_374, B[2], wc103);
  not gc103 (wc103, n_34);
  and g1895 (n_376, B[2], wc104);
  not gc104 (wc104, n_34);
  or g1896 (n_406, B[1], wc105);
  not gc105 (wc105, n_34);
  and g1897 (n_408, B[1], wc106);
  not gc106 (wc106, n_34);
  or g1898 (n_443, wc107, n_1783);
  not gc107 (wc107, n_34);
  and g1899 (n_445, wc108, n_1783);
  not gc108 (wc108, n_34);
  or g1900 (n_1824, n_376, wc109);
  not gc109 (wc109, n_374);
  or g1901 (n_1825, n_408, wc110);
  not gc110 (wc110, n_406);
  or g1902 (n_1826, n_445, wc111);
  not gc111 (wc111, n_443);
  or g1903 (n_1827, wc112, n_375);
  not gc112 (wc112, n_381);
  or g1904 (n_1828, wc113, n_407);
  not gc113 (wc113, n_413);
  or g1905 (n_1829, wc114, n_444);
  not gc114 (wc114, n_450);
  or g1906 (n_48, wc115, n_1751);
  not gc115 (wc115, n_1827);
  or g1907 (n_50, wc116, n_424);
  not gc116 (wc116, n_1828);
  or g1908 (n_1830, wc117, n_461);
  not gc117 (wc117, n_1829);
  and g1909 (n_51, n_50, wc118);
  not gc118 (wc118, n_48);
  or g1910 (n_53, n_1823, n_1830);
  and g1911 (n_54, n_53, wc119);
  not gc119 (wc119, n_50);
  or g1912 (n_58, wc120, wc121, wc122, wc123);
  and gc124 (wc123, wc124, n_47);
  not gc123 (wc124, n_53);
  and gc122 (wc122, n_54, n_46);
  and gc121 (wc121, n_51, n_45);
  and gc120 (wc120, n_48, n_34);
  or g1913 (n_56, wc125, wc126, wc128, wc129);
  and gc131 (wc129, wc130, wc131);
  not gc130 (wc131, n_1754);
  not gc129 (wc130, n_53);
  and gc128 (wc128, A[12], n_54);
  and gc127 (wc126, n_51, wc127);
  not gc126 (wc127, n_1754);
  and gc125 (wc125, A[12], n_48);
  or g1914 (n_57, wc132, wc133, wc134, wc135);
  and gc136 (wc135, wc136, n_44);
  not gc135 (wc136, n_53);
  and gc134 (wc134, n_54, n_1786);
  and gc133 (wc133, n_51, n_43);
  and gc132 (wc132, A[13], n_48);
  or g1915 (n_492, B[4], wc137);
  not gc137 (wc137, n_58);
  or g1916 (n_486, B[2], wc138);
  not gc138 (wc138, n_56);
  and g1917 (n_487, B[3], wc139);
  not gc139 (wc139, n_57);
  or g1918 (n_488, B[3], wc140);
  not gc140 (wc140, n_57);
  and g1919 (n_491, B[2], wc141);
  not gc141 (wc141, n_56);
  and g1920 (n_494, B[4], wc142);
  not gc142 (wc142, n_58);
  or g1921 (n_540, B[3], wc143);
  not gc143 (wc143, n_58);
  or g1922 (n_534, B[1], wc144);
  not gc144 (wc144, n_56);
  and g1923 (n_535, B[2], wc145);
  not gc145 (wc145, n_57);
  or g1924 (n_536, B[2], wc146);
  not gc146 (wc146, n_57);
  and g1925 (n_539, B[1], wc147);
  not gc147 (wc147, n_56);
  and g1926 (n_542, B[3], wc148);
  not gc148 (wc148, n_58);
  or g1927 (n_595, wc149, n_37);
  not gc149 (wc149, n_58);
  or g1928 (n_589, wc150, n_1783);
  not gc150 (wc150, n_56);
  and g1929 (n_590, wc151, n_36);
  not gc151 (wc151, n_57);
  or g1930 (n_591, wc152, n_36);
  not gc152 (wc152, n_57);
  and g1931 (n_594, wc153, n_1783);
  not gc153 (wc153, n_56);
  and g1932 (n_597, wc154, n_37);
  not gc154 (wc154, n_58);
  and g1933 (n_1831, n_488, wc155);
  not gc155 (wc155, n_489);
  or g1934 (n_1832, B[6], wc156);
  not gc156 (wc156, n_503);
  and g1935 (n_1833, n_536, wc157);
  not gc157 (wc157, n_537);
  and g1936 (n_1834, n_591, wc158);
  not gc158 (wc158, n_592);
  or g1937 (n_1835, n_494, wc159);
  not gc159 (wc159, n_492);
  or g1938 (n_1836, n_542, wc160);
  not gc160 (wc160, n_540);
  or g1939 (n_1837, n_597, wc161);
  not gc161 (wc161, n_595);
  or g1940 (n_1838, n_491, wc162);
  not gc162 (wc162, n_486);
  or g1941 (n_1839, n_539, wc163);
  not gc163 (wc163, n_534);
  or g1942 (n_1840, n_594, wc164);
  not gc164 (wc164, n_589);
  or g1943 (n_1841, n_491, wc165);
  not gc165 (wc165, n_495);
  or g1944 (n_1842, wc166, n_487);
  not gc166 (wc166, n_488);
  or g1945 (n_1843, n_539, wc167);
  not gc167 (wc167, n_543);
  or g1946 (n_1844, wc168, n_535);
  not gc168 (wc168, n_536);
  or g1947 (n_1845, n_594, wc169);
  not gc169 (wc169, n_598);
  or g1948 (n_1846, wc170, n_590);
  not gc170 (wc170, n_591);
  and g1949 (n_1847, wc171, n_493);
  not gc171 (wc171, B[6]);
  and g1950 (n_1848, n_310, n_541);
  and g1951 (n_1849, n_453, n_596);
  or g1952 (n_1850, n_1832, wc172);
  not gc172 (wc172, n_505);
  or g1953 (n_1851, n_563, wc173);
  not gc173 (wc173, n_556);
  or g1954 (n_1852, n_618, wc174);
  not gc174 (wc174, n_611);
  or g1955 (n_480, wc175, n_1847);
  not gc175 (wc175, n_1850);
  or g1956 (n_528, wc176, n_1848);
  not gc176 (wc176, n_1851);
  or g1957 (n_1853, wc177, n_1849);
  not gc177 (wc177, n_1852);
  or g1958 (n_74, wc178, n_1823);
  not gc178 (wc178, n_1853);
  and g1959 (n_73, wc179, n_480);
  not gc179 (wc179, n_528);
  or g1960 (n_81, wc180, wc182, wc183, wc184);
  and gc185 (wc184, wc185, n_70);
  not gc184 (wc185, n_74);
  and gc183 (wc183, n_69, n_75);
  and gc182 (wc182, n_73, n_68);
  and gc181 (wc180, wc181, n_58);
  not gc180 (wc181, n_480);
  or g1961 (n_79, wc186, wc188, wc189, wc190);
  and gc191 (wc190, wc191, n_64);
  not gc190 (wc191, n_74);
  and gc189 (wc189, n_63, n_75);
  and gc188 (wc188, n_73, n_62);
  and gc187 (wc186, wc187, n_56);
  not gc186 (wc187, n_480);
  or g1962 (n_80, wc192, wc194, wc195, wc196);
  and gc197 (wc196, wc197, n_67);
  not gc196 (wc197, n_74);
  and gc195 (wc195, n_66, n_75);
  and gc194 (wc194, n_73, n_65);
  and gc193 (wc192, wc193, n_57);
  not gc192 (wc193, n_480);
  or g1963 (n_77, wc198, wc200, wc202, wc203);
  and gc205 (wc203, wc204, wc205);
  not gc204 (wc205, n_1756);
  not gc203 (wc204, n_74);
  and gc202 (wc202, A[10], n_75);
  and gc201 (wc200, n_73, wc201);
  not gc200 (wc201, n_1756);
  and gc199 (wc198, A[10], wc199);
  not gc198 (wc199, n_480);
  or g1964 (n_78, wc206, wc208, wc209, wc210);
  and gc211 (wc210, wc211, n_61);
  not gc210 (wc211, n_74);
  and gc209 (wc209, n_1789, n_75);
  and gc208 (wc208, n_73, n_60);
  and gc207 (wc206, A[11], wc207);
  not gc206 (wc207, n_480);
  and g1965 (n_667, B[6], wc212);
  not gc212 (wc212, n_81);
  or g1966 (n_655, B[4], wc213);
  not gc213 (wc213, n_79);
  and g1967 (n_656, B[5], wc214);
  not gc214 (wc214, n_80);
  or g1968 (n_657, B[5], wc215);
  not gc215 (wc215, n_80);
  or g1969 (n_669, B[6], wc216);
  not gc216 (wc216, n_81);
  or g1970 (n_649, B[2], wc217);
  not gc217 (wc217, n_77);
  and g1971 (n_650, B[3], wc218);
  not gc218 (wc218, n_78);
  or g1972 (n_651, B[3], wc219);
  not gc219 (wc219, n_78);
  and g1973 (n_654, B[2], wc220);
  not gc220 (wc220, n_77);
  and g1974 (n_660, B[4], wc221);
  not gc221 (wc221, n_79);
  or g1975 (n_714, B[3], wc222);
  not gc222 (wc222, n_79);
  and g1976 (n_715, B[4], wc223);
  not gc223 (wc223, n_80);
  or g1977 (n_716, B[4], wc224);
  not gc224 (wc224, n_80);
  and g1978 (n_722, B[5], wc225);
  not gc225 (wc225, n_81);
  or g1979 (n_720, B[5], wc226);
  not gc226 (wc226, n_81);
  or g1980 (n_708, B[1], wc227);
  not gc227 (wc227, n_77);
  and g1981 (n_709, B[2], wc228);
  not gc228 (wc228, n_78);
  or g1982 (n_710, B[2], wc229);
  not gc229 (wc229, n_78);
  and g1983 (n_713, B[1], wc230);
  not gc230 (wc230, n_77);
  and g1984 (n_719, B[3], wc231);
  not gc231 (wc231, n_79);
  or g1985 (n_781, wc232, n_37);
  not gc232 (wc232, n_79);
  and g1986 (n_782, wc233, n_38);
  not gc233 (wc233, n_80);
  or g1987 (n_783, wc234, n_38);
  not gc234 (wc234, n_80);
  and g1988 (n_789, wc235, n_39);
  not gc235 (wc235, n_81);
  or g1989 (n_787, wc236, n_39);
  not gc236 (wc236, n_81);
  or g1990 (n_775, wc237, n_1783);
  not gc237 (wc237, n_77);
  and g1991 (n_776, wc238, n_36);
  not gc238 (wc238, n_78);
  or g1992 (n_777, wc239, n_36);
  not gc239 (wc239, n_78);
  and g1993 (n_780, wc240, n_1783);
  not gc240 (wc240, n_77);
  and g1994 (n_786, wc241, n_37);
  not gc241 (wc241, n_79);
  and g1995 (n_668, n_657, wc242);
  not gc242 (wc242, n_658);
  and g1996 (n_1854, n_651, wc243);
  not gc243 (wc243, n_652);
  or g1997 (n_1855, n_667, wc244);
  not gc244 (wc244, n_672);
  and g1998 (n_729, n_716, wc245);
  not gc245 (wc245, n_717);
  and g1999 (n_1856, n_710, wc246);
  not gc246 (wc246, n_711);
  and g2000 (n_796, n_783, wc247);
  not gc247 (wc247, n_784);
  and g2001 (n_1857, n_777, wc248);
  not gc248 (wc248, n_778);
  or g2002 (n_1858, wc249, n_667);
  not gc249 (wc249, n_669);
  or g2003 (n_1859, wc250, n_722);
  not gc250 (wc250, n_720);
  or g2004 (n_1860, wc251, n_789);
  not gc251 (wc251, n_787);
  or g2005 (n_1861, n_654, wc252);
  not gc252 (wc252, n_649);
  or g2006 (n_1862, n_713, wc253);
  not gc253 (wc253, n_708);
  or g2007 (n_1863, n_780, wc254);
  not gc254 (wc254, n_775);
  or g2008 (n_1864, n_654, wc255);
  not gc255 (wc255, n_661);
  or g2009 (n_1865, wc256, n_650);
  not gc256 (wc256, n_651);
  or g2010 (n_1866, n_713, wc257);
  not gc257 (wc257, n_723);
  or g2011 (n_1867, wc258, n_709);
  not gc258 (wc258, n_710);
  or g2012 (n_1868, n_780, wc259);
  not gc259 (wc259, n_790);
  or g2013 (n_1869, wc260, n_776);
  not gc260 (wc260, n_777);
  or g2014 (n_1870, n_660, wc261);
  not gc261 (wc261, n_655);
  or g2015 (n_1871, n_719, wc262);
  not gc262 (wc262, n_714);
  or g2016 (n_1872, n_786, wc263);
  not gc263 (wc263, n_781);
  or g2017 (n_1873, wc264, n_656);
  not gc264 (wc264, n_657);
  or g2018 (n_1874, wc265, n_715);
  not gc265 (wc265, n_716);
  or g2019 (n_1875, wc266, n_782);
  not gc266 (wc266, n_783);
  and g2020 (n_1876, wc267, n_734);
  not gc267 (wc267, n_729);
  and g2021 (n_1877, wc268, n_801);
  not gc268 (wc268, n_796);
  and g2022 (n_1878, n_669, wc269);
  not gc269 (wc269, n_670);
  or g2023 (n_1879, n_1855, wc270);
  not gc270 (wc270, n_674);
  or g2024 (n_1880, n_745, wc271);
  not gc271 (wc271, n_737);
  or g2025 (n_1881, n_812, wc272);
  not gc272 (wc272, n_804);
  or g2026 (n_1882, n_660, wc273);
  not gc273 (wc273, n_674);
  or g2027 (n_1883, n_719, wc274);
  not gc274 (wc274, n_737);
  or g2028 (n_1884, n_786, wc275);
  not gc275 (wc275, n_804);
  or g2029 (n_104, n_1823, wc276);
  not gc276 (wc276, n_816);
  and g2030 (n_102, wc277, n_643);
  not gc277 (wc277, n_702);
  or g2031 (n_116, wc278, wc280, wc281, wc282);
  and gc283 (wc282, wc283, n_99);
  not gc282 (wc283, n_104);
  and gc281 (wc281, n_98, n_105);
  and gc280 (wc280, n_102, n_97);
  and gc279 (wc278, n_81, wc279);
  not gc278 (wc279, n_643);
  or g2032 (n_112, wc284, wc286, wc287, wc288);
  and gc289 (wc288, wc289, n_87);
  not gc288 (wc289, n_104);
  and gc287 (wc287, n_86, n_105);
  and gc286 (wc286, n_102, n_85);
  and gc285 (wc284, n_77, wc285);
  not gc284 (wc285, n_643);
  or g2033 (n_113, wc290, wc292, wc293, wc294);
  and gc295 (wc294, wc295, n_90);
  not gc294 (wc295, n_104);
  and gc293 (wc293, n_89, n_105);
  and gc292 (wc292, n_102, n_88);
  and gc291 (wc290, n_78, wc291);
  not gc290 (wc291, n_643);
  or g2034 (n_114, wc296, wc298, wc299, wc300);
  and gc301 (wc300, wc301, n_93);
  not gc300 (wc301, n_104);
  and gc299 (wc299, n_92, n_105);
  and gc298 (wc298, n_102, n_91);
  and gc297 (wc296, n_79, wc297);
  not gc296 (wc297, n_643);
  or g2035 (n_115, wc302, wc304, wc305, wc306);
  and gc307 (wc306, wc307, n_96);
  not gc306 (wc307, n_104);
  and gc305 (wc305, n_95, n_105);
  and gc304 (wc304, n_102, n_94);
  and gc303 (wc302, n_80, wc303);
  not gc302 (wc303, n_643);
  or g2036 (n_110, wc308, wc310, wc312, wc313);
  and gc315 (wc313, wc314, wc315);
  not gc314 (wc315, n_1758);
  not gc313 (wc314, n_104);
  and gc312 (wc312, A[8], n_105);
  and gc311 (wc310, n_102, wc311);
  not gc310 (wc311, n_1758);
  and gc309 (wc308, A[8], wc309);
  not gc308 (wc309, n_643);
  or g2037 (n_111, wc316, wc318, wc319, wc320);
  and gc321 (wc320, wc321, n_84);
  not gc320 (wc321, n_104);
  and gc319 (wc319, n_1792, n_105);
  and gc318 (wc318, n_102, n_83);
  and gc317 (wc316, A[9], wc317);
  not gc316 (wc317, n_643);
  or g2038 (n_851, B[4], wc322);
  not gc322 (wc322, n_112);
  and g2039 (n_852, B[5], wc323);
  not gc323 (wc323, n_113);
  or g2040 (n_853, B[5], wc324);
  not gc324 (wc324, n_113);
  and g2041 (n_858, B[6], wc325);
  not gc325 (wc325, n_114);
  or g2042 (n_857, B[6], wc326);
  not gc326 (wc326, n_114);
  or g2043 (n_845, B[2], wc327);
  not gc327 (wc327, n_110);
  and g2044 (n_846, B[3], wc328);
  not gc328 (wc328, n_111);
  or g2045 (n_847, B[3], wc329);
  not gc329 (wc329, n_111);
  and g2046 (n_850, B[2], wc330);
  not gc330 (wc330, n_110);
  and g2047 (n_856, B[4], wc331);
  not gc331 (wc331, n_112);
  or g2048 (n_919, B[3], wc332);
  not gc332 (wc332, n_112);
  and g2049 (n_920, B[4], wc333);
  not gc333 (wc333, n_113);
  or g2050 (n_921, B[4], wc334);
  not gc334 (wc334, n_113);
  and g2051 (n_930, B[5], wc335);
  not gc335 (wc335, n_114);
  and g2052 (n_926, B[6], wc336);
  not gc336 (wc336, n_115);
  or g2053 (n_925, B[5], wc337);
  not gc337 (wc337, n_114);
  or g2054 (n_1885, B[6], wc338);
  not gc338 (wc338, n_115);
  or g2055 (n_913, B[1], wc339);
  not gc339 (wc339, n_110);
  and g2056 (n_914, B[2], wc340);
  not gc340 (wc340, n_111);
  or g2057 (n_915, B[2], wc341);
  not gc341 (wc341, n_111);
  and g2058 (n_918, B[1], wc342);
  not gc342 (wc342, n_110);
  and g2059 (n_924, B[3], wc343);
  not gc343 (wc343, n_112);
  or g2060 (n_1886, wc344, n_1823);
  not gc344 (wc344, n_116);
  or g2061 (n_999, wc345, n_37);
  not gc345 (wc345, n_112);
  and g2062 (n_1000, wc346, n_38);
  not gc346 (wc346, n_113);
  or g2063 (n_1001, wc347, n_38);
  not gc347 (wc347, n_113);
  and g2064 (n_1010, wc348, n_39);
  not gc348 (wc348, n_114);
  and g2065 (n_1006, wc349, n_40);
  not gc349 (wc349, n_115);
  or g2066 (n_1005, wc350, n_39);
  not gc350 (wc350, n_114);
  or g2067 (n_1887, wc351, n_40);
  not gc351 (wc351, n_115);
  or g2068 (n_993, wc352, n_1783);
  not gc352 (wc352, n_110);
  and g2069 (n_994, wc353, n_36);
  not gc353 (wc353, n_111);
  or g2070 (n_995, wc354, n_36);
  not gc354 (wc354, n_111);
  and g2071 (n_998, wc355, n_1783);
  not gc355 (wc355, n_110);
  and g2072 (n_1004, wc356, n_37);
  not gc356 (wc356, n_112);
  and g2073 (n_1888, wc357, n_1823);
  not gc357 (wc357, n_116);
  and g2074 (n_865, n_853, wc358);
  not gc358 (wc358, n_854);
  and g2075 (n_1889, n_857, wc359);
  not gc359 (wc359, n_115);
  and g2076 (n_1890, n_847, wc360);
  not gc360 (wc360, n_848);
  or g2077 (n_1891, n_858, wc361);
  not gc361 (wc361, n_868);
  and g2078 (n_937, n_921, wc362);
  not gc362 (wc362, n_922);
  and g2079 (n_1892, n_1885, wc363);
  not gc363 (wc363, n_928);
  and g2080 (n_1893, n_915, wc364);
  not gc364 (wc364, n_916);
  and g2081 (n_1017, n_1001, wc365);
  not gc365 (wc365, n_1002);
  and g2082 (n_1894, n_1887, wc366);
  not gc366 (wc366, n_1008);
  and g2083 (n_1895, n_995, wc367);
  not gc367 (wc367, n_996);
  or g2084 (n_1896, wc368, n_858);
  not gc368 (wc368, n_857);
  or g2085 (n_1897, wc369, n_930);
  not gc369 (wc369, n_925);
  or g2086 (n_1898, wc370, n_1010);
  not gc370 (wc370, n_1005);
  or g2087 (n_1899, n_850, wc371);
  not gc371 (wc371, n_845);
  or g2088 (n_1900, n_918, wc372);
  not gc372 (wc372, n_913);
  or g2089 (n_1901, n_998, wc373);
  not gc373 (wc373, n_993);
  or g2090 (n_1902, n_850, wc374);
  not gc374 (wc374, n_859);
  or g2091 (n_1903, wc375, n_846);
  not gc375 (wc375, n_847);
  or g2092 (n_1904, n_918, wc376);
  not gc376 (wc376, n_931);
  or g2093 (n_1905, wc377, n_914);
  not gc377 (wc377, n_915);
  or g2094 (n_1906, n_998, wc378);
  not gc378 (wc378, n_1011);
  or g2095 (n_1907, wc379, n_994);
  not gc379 (wc379, n_995);
  or g2096 (n_1908, n_856, wc380);
  not gc380 (wc380, n_851);
  or g2097 (n_1909, n_924, wc381);
  not gc381 (wc381, n_919);
  or g2098 (n_1910, n_1004, wc382);
  not gc382 (wc382, n_999);
  or g2099 (n_1911, wc383, n_852);
  not gc383 (wc383, n_853);
  or g2100 (n_1912, wc384, n_920);
  not gc384 (wc384, n_921);
  or g2101 (n_1913, wc385, n_1000);
  not gc385 (wc385, n_1001);
  and g2102 (n_1914, wc386, n_942);
  not gc386 (wc386, n_937);
  and g2103 (n_1915, wc387, n_1022);
  not gc387 (wc387, n_1017);
  and g2104 (n_1916, n_1889, wc388);
  not gc388 (wc388, n_871);
  or g2105 (n_1917, n_1891, wc389);
  not gc389 (wc389, n_873);
  and g2106 (n_1918, wc390, n_1892);
  not gc390 (wc390, n_1914);
  or g2107 (n_1919, n_955, wc391);
  not gc391 (wc391, n_947);
  and g2108 (n_1920, wc392, n_1894);
  not gc392 (wc392, n_1915);
  or g2109 (n_1921, n_1035, wc393);
  not gc393 (wc393, n_1027);
  or g2110 (n_1922, n_856, wc394);
  not gc394 (wc394, n_873);
  or g2111 (n_1923, n_924, wc395);
  not gc395 (wc395, n_947);
  or g2112 (n_1924, n_1004, wc396);
  not gc396 (wc396, n_1027);
  or g2113 (n_1925, n_1888, wc397);
  not gc397 (wc397, n_1040);
  or g2114 (n_839, n_882, n_116);
  or g2115 (n_907, n_959, n_116);
  and g2116 (n_147, wc398, n_839);
  not gc398 (wc398, n_907);
  and g2117 (n_150, n_907, wc399);
  not gc399 (wc399, n_151);
  or g2118 (n_161, wc400, wc402, wc403, wc404);
  and gc404 (wc404, n_137, n_151);
  and gc403 (wc403, n_150, n_136);
  and gc402 (wc402, n_147, n_135);
  and gc401 (wc400, wc401, n_114);
  not gc400 (wc401, n_839);
  or g2119 (n_157, wc405, wc407, wc408, wc409);
  and gc409 (wc409, n_125, n_151);
  and gc408 (wc408, n_150, n_124);
  and gc407 (wc407, n_147, n_123);
  and gc406 (wc405, wc406, n_110);
  not gc405 (wc406, n_839);
  or g2120 (n_158, wc410, wc412, wc413, wc414);
  and gc414 (wc414, n_128, n_151);
  and gc413 (wc413, n_150, n_127);
  and gc412 (wc412, n_147, n_126);
  and gc411 (wc410, wc411, n_111);
  not gc410 (wc411, n_839);
  or g2121 (n_159, wc415, wc417, wc418, wc419);
  and gc419 (wc419, n_131, n_151);
  and gc418 (wc418, n_150, n_130);
  and gc417 (wc417, n_147, n_129);
  and gc416 (wc415, wc416, n_112);
  not gc415 (wc416, n_839);
  or g2122 (n_160, wc420, wc422, wc423, wc424);
  and gc424 (wc424, n_134, n_151);
  and gc423 (wc423, n_150, n_133);
  and gc422 (wc422, n_147, n_132);
  and gc421 (wc420, wc421, n_113);
  not gc420 (wc421, n_839);
  or g2123 (n_155, wc425, wc427, wc429, wc430);
  and gc431 (wc430, wc431, n_151);
  not gc430 (wc431, n_1760);
  and gc429 (wc429, A[6], n_150);
  and gc428 (wc427, n_147, wc428);
  not gc427 (wc428, n_1760);
  and gc426 (wc425, A[6], wc426);
  not gc425 (wc426, n_839);
  or g2124 (n_156, wc432, wc434, wc435, wc436);
  and gc436 (wc436, n_122, n_151);
  and gc435 (wc435, n_150, n_1795);
  and gc434 (wc434, n_147, n_120);
  and gc433 (wc432, A[7], wc433);
  not gc432 (wc433, n_839);
  or g2125 (n_1080, B[4], wc437);
  not gc437 (wc437, n_157);
  and g2126 (n_1081, B[5], wc438);
  not gc438 (wc438, n_158);
  or g2127 (n_1082, B[5], wc439);
  not gc439 (wc439, n_158);
  and g2128 (n_1087, B[6], wc440);
  not gc440 (wc440, n_159);
  or g2129 (n_1086, B[6], wc441);
  not gc441 (wc441, n_159);
  or g2130 (n_1074, B[2], wc442);
  not gc442 (wc442, n_155);
  and g2131 (n_1075, B[3], wc443);
  not gc443 (wc443, n_156);
  or g2132 (n_1076, B[3], wc444);
  not gc444 (wc444, n_156);
  and g2133 (n_1079, B[2], wc445);
  not gc445 (wc445, n_155);
  and g2134 (n_1085, B[4], wc446);
  not gc446 (wc446, n_157);
  or g2135 (n_1148, B[3], wc447);
  not gc447 (wc447, n_157);
  and g2136 (n_1149, B[4], wc448);
  not gc448 (wc448, n_158);
  or g2137 (n_1150, B[4], wc449);
  not gc449 (wc449, n_158);
  and g2138 (n_1159, B[5], wc450);
  not gc450 (wc450, n_159);
  and g2139 (n_1155, B[6], wc451);
  not gc451 (wc451, n_160);
  or g2140 (n_1154, B[5], wc452);
  not gc452 (wc452, n_159);
  or g2141 (n_1926, B[6], wc453);
  not gc453 (wc453, n_160);
  or g2142 (n_1142, B[1], wc454);
  not gc454 (wc454, n_155);
  and g2143 (n_1143, B[2], wc455);
  not gc455 (wc455, n_156);
  or g2144 (n_1144, B[2], wc456);
  not gc456 (wc456, n_156);
  and g2145 (n_1147, B[1], wc457);
  not gc457 (wc457, n_155);
  and g2146 (n_1153, B[3], wc458);
  not gc458 (wc458, n_157);
  or g2147 (n_1927, wc459, n_1823);
  not gc459 (wc459, n_161);
  or g2148 (n_1228, wc460, n_37);
  not gc460 (wc460, n_157);
  and g2149 (n_1229, wc461, n_38);
  not gc461 (wc461, n_158);
  or g2150 (n_1230, wc462, n_38);
  not gc462 (wc462, n_158);
  and g2151 (n_1239, wc463, n_39);
  not gc463 (wc463, n_159);
  and g2152 (n_1235, wc464, n_40);
  not gc464 (wc464, n_160);
  or g2153 (n_1234, wc465, n_39);
  not gc465 (wc465, n_159);
  or g2154 (n_1928, wc466, n_40);
  not gc466 (wc466, n_160);
  or g2155 (n_1222, wc467, n_1783);
  not gc467 (wc467, n_155);
  and g2156 (n_1223, wc468, n_36);
  not gc468 (wc468, n_156);
  or g2157 (n_1224, wc469, n_36);
  not gc469 (wc469, n_156);
  and g2158 (n_1227, wc470, n_1783);
  not gc470 (wc470, n_155);
  and g2159 (n_1233, wc471, n_37);
  not gc471 (wc471, n_157);
  and g2160 (n_1929, wc472, n_1823);
  not gc472 (wc472, n_161);
  and g2161 (n_1094, n_1082, wc473);
  not gc473 (wc473, n_1083);
  and g2162 (n_1930, n_1086, wc474);
  not gc474 (wc474, n_160);
  and g2163 (n_1931, n_1076, wc475);
  not gc475 (wc475, n_1077);
  or g2164 (n_1932, n_1087, wc476);
  not gc476 (wc476, n_1097);
  and g2165 (n_1166, n_1150, wc477);
  not gc477 (wc477, n_1151);
  and g2166 (n_1933, n_1926, wc478);
  not gc478 (wc478, n_1157);
  and g2167 (n_1934, n_1144, wc479);
  not gc479 (wc479, n_1145);
  and g2168 (n_1246, n_1230, wc480);
  not gc480 (wc480, n_1231);
  and g2169 (n_1935, n_1928, wc481);
  not gc481 (wc481, n_1237);
  and g2170 (n_1936, n_1224, wc482);
  not gc482 (wc482, n_1225);
  or g2171 (n_1937, wc483, n_1087);
  not gc483 (wc483, n_1086);
  or g2172 (n_1938, wc484, n_1159);
  not gc484 (wc484, n_1154);
  or g2173 (n_1939, wc485, n_1239);
  not gc485 (wc485, n_1234);
  or g2174 (n_1940, n_1079, wc486);
  not gc486 (wc486, n_1074);
  or g2175 (n_1941, n_1147, wc487);
  not gc487 (wc487, n_1142);
  or g2176 (n_1942, n_1227, wc488);
  not gc488 (wc488, n_1222);
  or g2177 (n_1943, n_1079, wc489);
  not gc489 (wc489, n_1088);
  or g2178 (n_1944, wc490, n_1075);
  not gc490 (wc490, n_1076);
  or g2179 (n_1945, n_1147, wc491);
  not gc491 (wc491, n_1160);
  or g2180 (n_1946, wc492, n_1143);
  not gc492 (wc492, n_1144);
  or g2181 (n_1947, n_1227, wc493);
  not gc493 (wc493, n_1240);
  or g2182 (n_1948, wc494, n_1223);
  not gc494 (wc494, n_1224);
  or g2183 (n_1949, n_1085, wc495);
  not gc495 (wc495, n_1080);
  or g2184 (n_1950, n_1153, wc496);
  not gc496 (wc496, n_1148);
  or g2185 (n_1951, n_1233, wc497);
  not gc497 (wc497, n_1228);
  or g2186 (n_1952, wc498, n_1081);
  not gc498 (wc498, n_1082);
  or g2187 (n_1953, wc499, n_1149);
  not gc499 (wc499, n_1150);
  or g2188 (n_1954, wc500, n_1229);
  not gc500 (wc500, n_1230);
  and g2189 (n_1955, wc501, n_1171);
  not gc501 (wc501, n_1166);
  and g2190 (n_1956, wc502, n_1251);
  not gc502 (wc502, n_1246);
  and g2191 (n_1957, n_1930, wc503);
  not gc503 (wc503, n_1100);
  or g2192 (n_1958, n_1932, wc504);
  not gc504 (wc504, n_1102);
  and g2193 (n_1959, wc505, n_1933);
  not gc505 (wc505, n_1955);
  or g2194 (n_1960, n_1184, wc506);
  not gc506 (wc506, n_1176);
  and g2195 (n_1961, wc507, n_1935);
  not gc507 (wc507, n_1956);
  or g2196 (n_1962, n_1264, wc508);
  not gc508 (wc508, n_1256);
  or g2197 (n_1963, n_1085, wc509);
  not gc509 (wc509, n_1102);
  or g2198 (n_1964, n_1153, wc510);
  not gc510 (wc510, n_1176);
  or g2199 (n_1965, n_1233, wc511);
  not gc511 (wc511, n_1256);
  or g2200 (n_1966, n_1929, wc512);
  not gc512 (wc512, n_1269);
  or g2201 (n_1068, n_1111, n_161);
  or g2202 (n_1136, n_1188, n_161);
  and g2203 (n_192, wc513, n_1068);
  not gc513 (wc513, n_1136);
  and g2204 (n_195, n_1136, wc514);
  not gc514 (wc514, n_196);
  or g2205 (n_206, wc515, wc517, wc518, wc519);
  and gc519 (wc519, n_182, n_196);
  and gc518 (wc518, n_195, n_181);
  and gc517 (wc517, n_192, n_180);
  and gc516 (wc515, wc516, n_159);
  not gc515 (wc516, n_1068);
  or g2206 (n_202, wc520, wc522, wc523, wc524);
  and gc524 (wc524, n_170, n_196);
  and gc523 (wc523, n_195, n_169);
  and gc522 (wc522, n_192, n_168);
  and gc521 (wc520, wc521, n_155);
  not gc520 (wc521, n_1068);
  or g2207 (n_203, wc525, wc527, wc528, wc529);
  and gc529 (wc529, n_173, n_196);
  and gc528 (wc528, n_195, n_172);
  and gc527 (wc527, n_192, n_171);
  and gc526 (wc525, wc526, n_156);
  not gc525 (wc526, n_1068);
  or g2208 (n_204, wc530, wc532, wc533, wc534);
  and gc534 (wc534, n_176, n_196);
  and gc533 (wc533, n_195, n_175);
  and gc532 (wc532, n_192, n_174);
  and gc531 (wc530, wc531, n_157);
  not gc530 (wc531, n_1068);
  or g2209 (n_205, wc535, wc537, wc538, wc539);
  and gc539 (wc539, n_179, n_196);
  and gc538 (wc538, n_195, n_178);
  and gc537 (wc537, n_192, n_177);
  and gc536 (wc535, wc536, n_158);
  not gc535 (wc536, n_1068);
  or g2210 (n_200, wc540, wc542, wc544, wc545);
  and gc546 (wc545, wc546, n_196);
  not gc545 (wc546, n_1762);
  and gc544 (wc544, A[4], n_195);
  and gc543 (wc542, n_192, wc543);
  not gc542 (wc543, n_1762);
  and gc541 (wc540, A[4], wc541);
  not gc540 (wc541, n_1068);
  or g2211 (n_201, wc547, wc549, wc550, wc551);
  and gc551 (wc551, n_167, n_196);
  and gc550 (wc550, n_195, n_1798);
  and gc549 (wc549, n_192, n_165);
  and gc548 (wc547, A[5], wc548);
  not gc547 (wc548, n_1068);
  or g2212 (n_1309, B[4], wc552);
  not gc552 (wc552, n_202);
  and g2213 (n_1310, B[5], wc553);
  not gc553 (wc553, n_203);
  or g2214 (n_1311, B[5], wc554);
  not gc554 (wc554, n_203);
  and g2215 (n_1316, B[6], wc555);
  not gc555 (wc555, n_204);
  or g2216 (n_1315, B[6], wc556);
  not gc556 (wc556, n_204);
  or g2217 (n_1303, B[2], wc557);
  not gc557 (wc557, n_200);
  and g2218 (n_1304, B[3], wc558);
  not gc558 (wc558, n_201);
  or g2219 (n_1305, B[3], wc559);
  not gc559 (wc559, n_201);
  and g2220 (n_1308, B[2], wc560);
  not gc560 (wc560, n_200);
  and g2221 (n_1314, B[4], wc561);
  not gc561 (wc561, n_202);
  or g2222 (n_1377, B[3], wc562);
  not gc562 (wc562, n_202);
  and g2223 (n_1378, B[4], wc563);
  not gc563 (wc563, n_203);
  or g2224 (n_1379, B[4], wc564);
  not gc564 (wc564, n_203);
  and g2225 (n_1388, B[5], wc565);
  not gc565 (wc565, n_204);
  and g2226 (n_1384, B[6], wc566);
  not gc566 (wc566, n_205);
  or g2227 (n_1383, B[5], wc567);
  not gc567 (wc567, n_204);
  or g2228 (n_1967, B[6], wc568);
  not gc568 (wc568, n_205);
  or g2229 (n_1371, B[1], wc569);
  not gc569 (wc569, n_200);
  and g2230 (n_1372, B[2], wc570);
  not gc570 (wc570, n_201);
  or g2231 (n_1373, B[2], wc571);
  not gc571 (wc571, n_201);
  and g2232 (n_1376, B[1], wc572);
  not gc572 (wc572, n_200);
  and g2233 (n_1382, B[3], wc573);
  not gc573 (wc573, n_202);
  or g2234 (n_1968, wc574, n_1823);
  not gc574 (wc574, n_206);
  or g2235 (n_1457, wc575, n_37);
  not gc575 (wc575, n_202);
  and g2236 (n_1458, wc576, n_38);
  not gc576 (wc576, n_203);
  or g2237 (n_1459, wc577, n_38);
  not gc577 (wc577, n_203);
  and g2238 (n_1468, wc578, n_39);
  not gc578 (wc578, n_204);
  and g2239 (n_1464, wc579, n_40);
  not gc579 (wc579, n_205);
  or g2240 (n_1463, wc580, n_39);
  not gc580 (wc580, n_204);
  or g2241 (n_1969, wc581, n_40);
  not gc581 (wc581, n_205);
  or g2242 (n_1451, wc582, n_1783);
  not gc582 (wc582, n_200);
  and g2243 (n_1452, wc583, n_36);
  not gc583 (wc583, n_201);
  or g2244 (n_1453, wc584, n_36);
  not gc584 (wc584, n_201);
  and g2245 (n_1456, wc585, n_1783);
  not gc585 (wc585, n_200);
  and g2246 (n_1462, wc586, n_37);
  not gc586 (wc586, n_202);
  and g2247 (n_1970, wc587, n_1823);
  not gc587 (wc587, n_206);
  and g2248 (n_1323, n_1311, wc588);
  not gc588 (wc588, n_1312);
  and g2249 (n_1971, n_1315, wc589);
  not gc589 (wc589, n_205);
  and g2250 (n_1972, n_1305, wc590);
  not gc590 (wc590, n_1306);
  or g2251 (n_1973, n_1316, wc591);
  not gc591 (wc591, n_1326);
  and g2252 (n_1395, n_1379, wc592);
  not gc592 (wc592, n_1380);
  and g2253 (n_1974, n_1967, wc593);
  not gc593 (wc593, n_1386);
  and g2254 (n_1975, n_1373, wc594);
  not gc594 (wc594, n_1374);
  and g2255 (n_1475, n_1459, wc595);
  not gc595 (wc595, n_1460);
  and g2256 (n_1976, n_1969, wc596);
  not gc596 (wc596, n_1466);
  and g2257 (n_1977, n_1453, wc597);
  not gc597 (wc597, n_1454);
  or g2258 (n_1978, wc598, n_1316);
  not gc598 (wc598, n_1315);
  or g2259 (n_1979, wc599, n_1388);
  not gc599 (wc599, n_1383);
  or g2260 (n_1980, wc600, n_1468);
  not gc600 (wc600, n_1463);
  or g2261 (n_1981, n_1308, wc601);
  not gc601 (wc601, n_1303);
  or g2262 (n_1982, n_1376, wc602);
  not gc602 (wc602, n_1371);
  or g2263 (n_1983, n_1456, wc603);
  not gc603 (wc603, n_1451);
  or g2264 (n_1984, n_1308, wc604);
  not gc604 (wc604, n_1317);
  or g2265 (n_1985, wc605, n_1304);
  not gc605 (wc605, n_1305);
  or g2266 (n_1986, n_1376, wc606);
  not gc606 (wc606, n_1389);
  or g2267 (n_1987, wc607, n_1372);
  not gc607 (wc607, n_1373);
  or g2268 (n_1988, n_1456, wc608);
  not gc608 (wc608, n_1469);
  or g2269 (n_1989, wc609, n_1452);
  not gc609 (wc609, n_1453);
  or g2270 (n_1990, n_1314, wc610);
  not gc610 (wc610, n_1309);
  or g2271 (n_1991, n_1382, wc611);
  not gc611 (wc611, n_1377);
  or g2272 (n_1992, n_1462, wc612);
  not gc612 (wc612, n_1457);
  or g2273 (n_1993, wc613, n_1310);
  not gc613 (wc613, n_1311);
  or g2274 (n_1994, wc614, n_1378);
  not gc614 (wc614, n_1379);
  or g2275 (n_1995, wc615, n_1458);
  not gc615 (wc615, n_1459);
  and g2276 (n_1996, wc616, n_1400);
  not gc616 (wc616, n_1395);
  and g2277 (n_1997, wc617, n_1480);
  not gc617 (wc617, n_1475);
  and g2278 (n_1998, n_1971, wc618);
  not gc618 (wc618, n_1329);
  or g2279 (n_1999, n_1973, wc619);
  not gc619 (wc619, n_1331);
  and g2280 (n_2000, wc620, n_1974);
  not gc620 (wc620, n_1996);
  or g2281 (n_2001, n_1413, wc621);
  not gc621 (wc621, n_1405);
  and g2282 (n_2002, wc622, n_1976);
  not gc622 (wc622, n_1997);
  or g2283 (n_2003, n_1493, wc623);
  not gc623 (wc623, n_1485);
  or g2284 (n_2004, n_1314, wc624);
  not gc624 (wc624, n_1331);
  or g2285 (n_2005, n_1382, wc625);
  not gc625 (wc625, n_1405);
  or g2286 (n_2006, n_1462, wc626);
  not gc626 (wc626, n_1485);
  or g2287 (n_2007, n_1970, wc627);
  not gc627 (wc627, n_1498);
  or g2288 (n_1297, n_1340, n_206);
  or g2289 (n_1365, n_1417, n_206);
  and g2290 (n_237, wc628, n_1297);
  not gc628 (wc628, n_1365);
  and g2291 (n_240, n_1365, wc629);
  not gc629 (wc629, n_241);
  or g2292 (n_251, wc630, wc632, wc633, wc634);
  and gc634 (wc634, n_227, n_241);
  and gc633 (wc633, n_240, n_226);
  and gc632 (wc632, n_237, n_225);
  and gc631 (wc630, wc631, n_204);
  not gc630 (wc631, n_1297);
  or g2293 (n_247, wc635, wc637, wc638, wc639);
  and gc639 (wc639, n_215, n_241);
  and gc638 (wc638, n_240, n_214);
  and gc637 (wc637, n_237, n_213);
  and gc636 (wc635, wc636, n_200);
  not gc635 (wc636, n_1297);
  or g2294 (n_248, wc640, wc642, wc643, wc644);
  and gc644 (wc644, n_218, n_241);
  and gc643 (wc643, n_240, n_217);
  and gc642 (wc642, n_237, n_216);
  and gc641 (wc640, wc641, n_201);
  not gc640 (wc641, n_1297);
  or g2295 (n_249, wc645, wc647, wc648, wc649);
  and gc649 (wc649, n_221, n_241);
  and gc648 (wc648, n_240, n_220);
  and gc647 (wc647, n_237, n_219);
  and gc646 (wc645, wc646, n_202);
  not gc645 (wc646, n_1297);
  or g2296 (n_250, wc650, wc652, wc653, wc654);
  and gc654 (wc654, n_224, n_241);
  and gc653 (wc653, n_240, n_223);
  and gc652 (wc652, n_237, n_222);
  and gc651 (wc650, wc651, n_203);
  not gc650 (wc651, n_1297);
  or g2297 (n_245, wc655, wc657, wc659, wc660);
  and gc661 (wc660, wc661, n_241);
  not gc660 (wc661, n_1764);
  and gc659 (wc659, A[2], n_240);
  and gc658 (wc657, n_237, wc658);
  not gc657 (wc658, n_1764);
  and gc656 (wc655, A[2], wc656);
  not gc655 (wc656, n_1297);
  or g2298 (n_246, wc662, wc664, wc665, wc666);
  and gc666 (wc666, n_212, n_241);
  and gc665 (wc665, n_240, n_1801);
  and gc664 (wc664, n_237, n_210);
  and gc663 (wc662, A[3], wc663);
  not gc662 (wc663, n_1297);
  or g2299 (n_1538, B[4], wc667);
  not gc667 (wc667, n_247);
  and g2300 (n_1539, B[5], wc668);
  not gc668 (wc668, n_248);
  or g2301 (n_1540, B[5], wc669);
  not gc669 (wc669, n_248);
  and g2302 (n_1545, B[6], wc670);
  not gc670 (wc670, n_249);
  or g2303 (n_1544, B[6], wc671);
  not gc671 (wc671, n_249);
  or g2304 (n_1532, B[2], wc672);
  not gc672 (wc672, n_245);
  and g2305 (n_1533, B[3], wc673);
  not gc673 (wc673, n_246);
  or g2306 (n_1534, B[3], wc674);
  not gc674 (wc674, n_246);
  and g2307 (n_1537, B[2], wc675);
  not gc675 (wc675, n_245);
  and g2308 (n_1543, B[4], wc676);
  not gc676 (wc676, n_247);
  or g2309 (n_1606, B[3], wc677);
  not gc677 (wc677, n_247);
  and g2310 (n_1607, B[4], wc678);
  not gc678 (wc678, n_248);
  or g2311 (n_1608, B[4], wc679);
  not gc679 (wc679, n_248);
  and g2312 (n_1617, B[5], wc680);
  not gc680 (wc680, n_249);
  and g2313 (n_1613, B[6], wc681);
  not gc681 (wc681, n_250);
  or g2314 (n_1612, B[5], wc682);
  not gc682 (wc682, n_249);
  or g2315 (n_2008, B[6], wc683);
  not gc683 (wc683, n_250);
  or g2316 (n_1600, B[1], wc684);
  not gc684 (wc684, n_245);
  and g2317 (n_1601, B[2], wc685);
  not gc685 (wc685, n_246);
  or g2318 (n_1602, B[2], wc686);
  not gc686 (wc686, n_246);
  and g2319 (n_1605, B[1], wc687);
  not gc687 (wc687, n_245);
  and g2320 (n_1611, B[3], wc688);
  not gc688 (wc688, n_247);
  or g2321 (n_2009, wc689, n_1823);
  not gc689 (wc689, n_251);
  or g2322 (n_1686, wc690, n_37);
  not gc690 (wc690, n_247);
  and g2323 (n_1687, wc691, n_38);
  not gc691 (wc691, n_248);
  or g2324 (n_1688, wc692, n_38);
  not gc692 (wc692, n_248);
  and g2325 (n_1697, wc693, n_39);
  not gc693 (wc693, n_249);
  and g2326 (n_1693, wc694, n_40);
  not gc694 (wc694, n_250);
  or g2327 (n_1692, wc695, n_39);
  not gc695 (wc695, n_249);
  or g2328 (n_2010, wc696, n_40);
  not gc696 (wc696, n_250);
  or g2329 (n_1680, wc697, n_1783);
  not gc697 (wc697, n_245);
  and g2330 (n_1681, wc698, n_36);
  not gc698 (wc698, n_246);
  or g2331 (n_1682, wc699, n_36);
  not gc699 (wc699, n_246);
  and g2332 (n_1685, wc700, n_1783);
  not gc700 (wc700, n_245);
  and g2333 (n_1691, wc701, n_37);
  not gc701 (wc701, n_247);
  and g2334 (n_2011, wc702, n_1823);
  not gc702 (wc702, n_251);
  and g2335 (n_1552, n_1540, wc703);
  not gc703 (wc703, n_1541);
  and g2336 (n_2012, n_1544, wc704);
  not gc704 (wc704, n_250);
  and g2337 (n_2013, n_1534, wc705);
  not gc705 (wc705, n_1535);
  or g2338 (n_2014, n_1545, wc706);
  not gc706 (wc706, n_1555);
  and g2339 (n_1624, n_1608, wc707);
  not gc707 (wc707, n_1609);
  and g2340 (n_2015, n_2008, wc708);
  not gc708 (wc708, n_1615);
  and g2341 (n_2016, n_1602, wc709);
  not gc709 (wc709, n_1603);
  and g2342 (n_1704, n_1688, wc710);
  not gc710 (wc710, n_1689);
  and g2343 (n_2017, n_2010, wc711);
  not gc711 (wc711, n_1695);
  and g2344 (n_2018, n_1682, wc712);
  not gc712 (wc712, n_1683);
  or g2345 (n_2019, n_1537, wc713);
  not gc713 (wc713, n_1546);
  or g2346 (n_2020, n_1537, wc714);
  not gc714 (wc714, n_1532);
  or g2347 (n_2021, wc715, n_1533);
  not gc715 (wc715, n_1534);
  or g2348 (n_2022, n_1543, wc716);
  not gc716 (wc716, n_1538);
  or g2349 (n_2023, wc717, n_1539);
  not gc717 (wc717, n_1540);
  or g2350 (n_2024, wc718, n_1545);
  not gc718 (wc718, n_1544);
  or g2351 (n_2025, n_1605, wc719);
  not gc719 (wc719, n_1618);
  or g2352 (n_2026, n_1605, wc720);
  not gc720 (wc720, n_1600);
  or g2353 (n_2027, wc721, n_1601);
  not gc721 (wc721, n_1602);
  or g2354 (n_2028, n_1611, wc722);
  not gc722 (wc722, n_1606);
  or g2355 (n_2029, wc723, n_1607);
  not gc723 (wc723, n_1608);
  or g2356 (n_2030, wc724, n_1617);
  not gc724 (wc724, n_1612);
  or g2357 (n_2031, n_1685, wc725);
  not gc725 (wc725, n_1698);
  or g2358 (n_2032, n_1685, wc726);
  not gc726 (wc726, n_1680);
  or g2359 (n_2033, wc727, n_1681);
  not gc727 (wc727, n_1682);
  or g2360 (n_2034, n_1691, wc728);
  not gc728 (wc728, n_1686);
  or g2361 (n_2035, wc729, n_1687);
  not gc729 (wc729, n_1688);
  or g2362 (n_2036, wc730, n_1697);
  not gc730 (wc730, n_1692);
  and g2363 (n_2037, wc731, n_1629);
  not gc731 (wc731, n_1624);
  and g2364 (n_2038, wc732, n_1709);
  not gc732 (wc732, n_1704);
  and g2365 (n_2039, n_2012, wc733);
  not gc733 (wc733, n_1558);
  or g2366 (n_2040, n_2014, wc734);
  not gc734 (wc734, n_1560);
  and g2367 (n_2041, wc735, n_2015);
  not gc735 (wc735, n_2037);
  or g2368 (n_2042, n_1642, wc736);
  not gc736 (wc736, n_1634);
  and g2369 (n_2043, wc737, n_2017);
  not gc737 (wc737, n_2038);
  or g2370 (n_2044, n_1722, wc738);
  not gc738 (wc738, n_1714);
  or g2371 (n_2045, n_1543, wc739);
  not gc739 (wc739, n_1560);
  or g2372 (n_2046, n_1611, wc740);
  not gc740 (wc740, n_1634);
  or g2373 (n_2047, n_1691, wc741);
  not gc741 (wc741, n_1714);
  or g2374 (n_2048, n_2011, wc742);
  not gc742 (wc742, n_1727);
  or g2375 (n_1526, n_1569, n_251);
  or g2376 (n_1594, n_1646, n_251);
  and g2377 (n_282, wc743, n_1526);
  not gc743 (wc743, n_1594);
  and g2378 (n_285, n_1594, wc744);
  not gc744 (wc744, n_286);
  or g2379 (REMAINDER[6], wc745, wc747, wc748, wc749);
  and gc749 (wc749, n_272, n_286);
  and gc748 (wc748, n_285, n_271);
  and gc747 (wc747, n_282, n_270);
  and gc746 (wc745, wc746, n_249);
  not gc745 (wc746, n_1526);
  or g2380 (REMAINDER[5], wc750, wc752, wc753, wc754);
  and gc754 (wc754, n_269, n_286);
  and gc753 (wc753, n_285, n_268);
  and gc752 (wc752, n_282, n_267);
  and gc751 (wc750, wc751, n_248);
  not gc750 (wc751, n_1526);
  or g2381 (REMAINDER[4], wc755, wc757, wc758, wc759);
  and gc759 (wc759, n_266, n_286);
  and gc758 (wc758, n_285, n_265);
  and gc757 (wc757, n_282, n_264);
  and gc756 (wc755, wc756, n_247);
  not gc755 (wc756, n_1526);
  or g2382 (REMAINDER[3], wc760, wc762, wc763, wc764);
  and gc764 (wc764, n_263, n_286);
  and gc763 (wc763, n_285, n_262);
  and gc762 (wc762, n_282, n_261);
  and gc761 (wc760, wc761, n_246);
  not gc760 (wc761, n_1526);
  or g2383 (REMAINDER[2], wc765, wc767, wc768, wc769);
  and gc769 (wc769, n_260, n_286);
  and gc768 (wc768, n_285, n_259);
  and gc767 (wc767, n_282, n_258);
  and gc766 (wc765, wc766, n_245);
  not gc765 (wc766, n_1526);
  or g2384 (REMAINDER[1], wc770, wc772, wc773, wc774);
  and gc774 (wc774, n_257, n_286);
  and gc773 (wc773, n_285, n_1804);
  and gc772 (wc772, n_282, n_255);
  and gc771 (wc770, A[1], wc771);
  not gc770 (wc771, n_1526);
  or g2385 (REMAINDER[0], wc775, wc777, wc779, wc780);
  and gc781 (wc780, wc781, n_286);
  not gc780 (wc781, n_1766);
  and gc779 (wc779, A[0], n_285);
  and gc778 (wc777, n_282, wc778);
  not gc777 (wc778, n_1766);
  and gc776 (wc775, A[0], wc776);
  not gc775 (wc776, n_1526);
endmodule

module remainder_unsigned_GENERIC(A, B, REMAINDER);
  input [14:0] A;
  input [6:0] B;
  output [14:0] REMAINDER;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] REMAINDER;
  remainder_unsigned_GENERIC_REAL g1(.A (A), .B (B), .REMAINDER
       (REMAINDER));
endmodule

module remainder_unsigned_268_GENERIC_REAL(A, B, REMAINDER);
// synthesis_equation "assign REMAINDER = A % B;"
  input [14:0] A;
  input [6:0] B;
  output [14:0] REMAINDER;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] REMAINDER;
  wire n_32, n_34, n_36, n_37, n_38, n_39, n_40, n_43;
  wire n_44, n_45, n_46, n_47, n_48, n_50, n_51, n_53;
  wire n_54, n_56, n_57, n_58, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_73;
  wire n_74, n_75, n_77, n_78, n_79, n_80, n_81, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_102, n_104, n_105, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_120, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_147, n_150, n_151, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_165, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_192, n_195;
  wire n_196, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_210, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_237, n_240, n_241, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_255, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_282, n_285, n_286, n_295;
  wire n_298, n_301, n_303, n_304, n_305, n_306, n_309, n_310;
  wire n_311, n_312, n_315, n_318, n_320, n_322, n_324, n_325;
  wire n_328, n_329, n_335, n_339, n_341, n_342, n_351, n_353;
  wire n_370, n_372, n_374, n_375, n_376, n_377, n_380, n_381;
  wire n_401, n_404, n_406, n_407, n_408, n_409, n_412, n_413;
  wire n_424, n_441, n_443, n_444, n_445, n_446, n_449, n_450;
  wire n_451, n_453, n_461, n_480, n_482, n_484, n_486, n_487;
  wire n_488, n_489, n_491, n_492, n_493, n_494, n_495, n_498;
  wire n_500, n_503, n_505, n_515, n_528, n_529, n_532, n_534;
  wire n_535, n_536, n_537, n_539, n_540, n_541, n_542, n_543;
  wire n_546, n_548, n_551, n_556, n_563, n_569, n_587, n_589;
  wire n_590, n_591, n_592, n_594, n_595, n_596, n_597, n_598;
  wire n_601, n_603, n_606, n_611, n_618, n_626, n_643, n_645;
  wire n_647, n_649, n_650, n_651, n_652, n_654, n_655, n_656;
  wire n_657, n_658, n_660, n_661, n_664, n_666, n_667, n_668;
  wire n_669, n_670, n_672, n_674, n_677, n_685, n_689, n_691;
  wire n_702, n_703, n_706, n_708, n_709, n_710, n_711, n_713;
  wire n_714, n_715, n_716, n_717, n_719, n_720, n_721, n_722;
  wire n_723, n_726, n_728, n_729, n_732, n_734, n_737, n_740;
  wire n_745, n_747, n_752, n_756, n_758, n_773, n_775, n_776;
  wire n_777, n_778, n_780, n_781, n_782, n_783, n_784, n_786;
  wire n_787, n_788, n_789, n_790, n_793, n_795, n_796, n_799;
  wire n_801, n_804, n_807, n_812, n_814, n_816, n_821, n_825;
  wire n_827, n_839, n_841, n_843, n_845, n_846, n_847, n_848;
  wire n_850, n_851, n_852, n_853, n_854, n_856, n_857, n_858;
  wire n_859, n_862, n_864, n_865, n_868, n_871, n_873, n_876;
  wire n_882, n_887, n_891, n_893, n_907, n_908, n_911, n_913;
  wire n_914, n_915, n_916, n_918, n_919, n_920, n_921, n_922;
  wire n_924, n_925, n_926, n_928, n_930, n_931, n_934, n_936;
  wire n_937, n_940, n_942, n_947, n_950, n_955, n_959, n_964;
  wire n_968, n_970, n_991, n_993, n_994, n_995, n_996, n_998;
  wire n_999, n_1000, n_1001, n_1002, n_1004, n_1005, n_1006, n_1008;
  wire n_1010, n_1011, n_1014, n_1016, n_1017, n_1020, n_1022, n_1027;
  wire n_1030, n_1035, n_1040, n_1047, n_1051, n_1053, n_1068, n_1070;
  wire n_1072, n_1074, n_1075, n_1076, n_1077, n_1079, n_1080, n_1081;
  wire n_1082, n_1083, n_1085, n_1086, n_1087, n_1088, n_1091, n_1093;
  wire n_1094, n_1097, n_1100, n_1102, n_1105, n_1111, n_1116, n_1120;
  wire n_1122, n_1136, n_1137, n_1140, n_1142, n_1143, n_1144, n_1145;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1153, n_1154, n_1155;
  wire n_1157, n_1159, n_1160, n_1163, n_1165, n_1166, n_1169, n_1171;
  wire n_1176, n_1179, n_1184, n_1188, n_1193, n_1197, n_1199, n_1220;
  wire n_1222, n_1223, n_1224, n_1225, n_1227, n_1228, n_1229, n_1230;
  wire n_1231, n_1233, n_1234, n_1235, n_1237, n_1239, n_1240, n_1243;
  wire n_1245, n_1246, n_1249, n_1251, n_1256, n_1259, n_1264, n_1269;
  wire n_1276, n_1280, n_1282, n_1297, n_1299, n_1301, n_1303, n_1304;
  wire n_1305, n_1306, n_1308, n_1309, n_1310, n_1311, n_1312, n_1314;
  wire n_1315, n_1316, n_1317, n_1320, n_1322, n_1323, n_1326, n_1329;
  wire n_1331, n_1334, n_1340, n_1345, n_1349, n_1351, n_1365, n_1366;
  wire n_1369, n_1371, n_1372, n_1373, n_1374, n_1376, n_1377, n_1378;
  wire n_1379, n_1380, n_1382, n_1383, n_1384, n_1386, n_1388, n_1389;
  wire n_1392, n_1394, n_1395, n_1398, n_1400, n_1405, n_1408, n_1413;
  wire n_1417, n_1422, n_1426, n_1428, n_1449, n_1451, n_1452, n_1453;
  wire n_1454, n_1456, n_1457, n_1458, n_1459, n_1460, n_1462, n_1463;
  wire n_1464, n_1466, n_1468, n_1469, n_1472, n_1474, n_1475, n_1478;
  wire n_1480, n_1485, n_1488, n_1493, n_1498, n_1505, n_1509, n_1511;
  wire n_1526, n_1528, n_1530, n_1532, n_1533, n_1534, n_1535, n_1537;
  wire n_1538, n_1539, n_1540, n_1541, n_1543, n_1544, n_1545, n_1546;
  wire n_1549, n_1551, n_1552, n_1555, n_1558, n_1560, n_1563, n_1569;
  wire n_1574, n_1578, n_1580, n_1594, n_1595, n_1598, n_1600, n_1601;
  wire n_1602, n_1603, n_1605, n_1606, n_1607, n_1608, n_1609, n_1611;
  wire n_1612, n_1613, n_1615, n_1617, n_1618, n_1621, n_1623, n_1624;
  wire n_1627, n_1629, n_1634, n_1637, n_1642, n_1646, n_1651, n_1655;
  wire n_1657, n_1678, n_1680, n_1681, n_1682, n_1683, n_1685, n_1686;
  wire n_1687, n_1688, n_1689, n_1691, n_1692, n_1693, n_1695, n_1697;
  wire n_1698, n_1701, n_1703, n_1704, n_1707, n_1709, n_1714, n_1717;
  wire n_1722, n_1727, n_1734, n_1738, n_1740, n_1750, n_1751, n_1752;
  wire n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760;
  wire n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768;
  wire n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832;
  wire n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840;
  wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864;
  wire n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872;
  wire n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880;
  wire n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888;
  wire n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896;
  wire n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904;
  wire n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912;
  wire n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920;
  wire n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928;
  wire n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936;
  wire n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960;
  wire n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976;
  wire n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984;
  wire n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992;
  wire n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000;
  wire n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016;
  wire n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024;
  wire n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032;
  wire n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040;
  wire n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048;
  assign REMAINDER[7] = 1'b0;
  assign REMAINDER[8] = 1'b0;
  assign REMAINDER[9] = 1'b0;
  assign REMAINDER[10] = 1'b0;
  assign REMAINDER[11] = 1'b0;
  assign REMAINDER[12] = 1'b0;
  assign REMAINDER[13] = 1'b0;
  assign REMAINDER[14] = 1'b0;
  and g19 (n_75, n_528, n_74);
  and g31 (n_105, n_702, n_104);
  xor g84 (n_342, B[0], B[1]);
  nand g2 (n_295, B[0], B[1]);
  nor g87 (n_298, B[1], B[2]);
  nand g88 (n_301, B[1], B[2]);
  nand g90 (n_303, B[2], B[3]);
  nand g92 (n_305, B[3], B[4]);
  nand g13 (n_309, B[4], B[5]);
  nand g15 (n_311, B[5], B[6]);
  nand g95 (n_315, n_301, n_1769);
  nor g96 (n_306, n_303, n_304);
  nor g24 (n_318, n_351, n_304);
  nor g25 (n_312, n_309, n_310);
  nor g99 (n_324, n_353, n_310);
  nand g102 (n_335, n_303, n_1807);
  nand g103 (n_320, n_318, n_315);
  nand g104 (n_325, n_1773, n_320);
  nand g38 (n_329, n_324, B[6]);
  nand g107 (n_339, n_309, n_1821);
  nand g108 (n_328, n_324, n_325);
  nand g109 (n_341, n_322, n_328);
  xnor g50 (n_36, n_315, n_1770);
  xnor g115 (n_37, n_335, n_1772);
  xnor g117 (n_38, n_325, n_1774);
  xnor g120 (n_39, n_339, n_1775);
  nor g126 (n_351, B[2], B[3]);
  nor g36 (n_353, B[4], B[5]);
  nand g158 (n_377, n_372, n_1782);
  nor g159 (n_375, n_374, B[3]);
  nor g160 (n_380, n_376, B[3]);
  nand g165 (n_381, n_380, n_377);
  xnor g175 (n_43, n_370, n_1785);
  xnor g177 (n_45, n_377, n_1824);
  nand g197 (n_409, n_404, n_401);
  nor g198 (n_407, n_406, B[2]);
  nor g199 (n_412, n_408, B[2]);
  nor g200 (n_304, B[3], B[4]);
  nor g201 (n_310, B[5], B[6]);
  nand g205 (n_413, n_412, n_409);
  nand g209 (n_424, n_304, n_310);
  xnor g220 (n_46, n_409, n_1825);
  nand g243 (n_446, n_441, n_1806);
  nor g244 (n_444, n_443, n_36);
  nor g245 (n_449, n_445, n_36);
  nor g246 (n_451, n_37, n_38);
  nor g247 (n_453, n_39, n_40);
  nand g251 (n_450, n_449, n_446);
  nand g255 (n_461, n_451, n_453);
  xnor g266 (n_44, n_370, n_1808);
  xnor g268 (n_47, n_446, n_1826);
  nand g303 (n_495, n_484, n_1787);
  nor g304 (n_489, n_486, n_487);
  nor g307 (n_498, n_491, n_487);
  nor g308 (n_493, n_492, B[5]);
  nor g309 (n_503, n_494, B[5]);
  nand g312 (n_515, n_486, n_1841);
  nand g313 (n_500, n_498, n_495);
  nand g314 (n_505, n_1831, n_500);
  xnor g327 (n_60, n_482, n_1788);
  xnor g329 (n_62, n_495, n_1838);
  xnor g332 (n_65, n_515, n_1842);
  xnor g334 (n_68, n_505, n_1835);
  nand g359 (n_543, n_532, n_529);
  nor g360 (n_537, n_534, n_535);
  nor g363 (n_546, n_539, n_535);
  nor g364 (n_541, n_540, B[4]);
  nor g365 (n_551, n_542, B[4]);
  nand g369 (n_569, n_534, n_1843);
  nand g370 (n_548, n_546, n_543);
  nand g371 (n_556, n_1833, n_548);
  nand g377 (n_563, n_551, n_310);
  xnor g392 (n_63, n_543, n_1839);
  xnor g395 (n_66, n_569, n_1844);
  xnor g397 (n_69, n_556, n_1836);
  nand g423 (n_598, n_587, n_1809);
  nor g424 (n_592, n_589, n_590);
  nor g427 (n_601, n_594, n_590);
  nor g428 (n_596, n_595, n_38);
  nor g429 (n_606, n_597, n_38);
  nand g433 (n_626, n_589, n_1845);
  nand g434 (n_603, n_601, n_598);
  nand g435 (n_611, n_1834, n_603);
  nand g441 (n_618, n_606, n_453);
  xnor g456 (n_61, n_482, n_1810);
  xnor g458 (n_64, n_598, n_1840);
  xnor g461 (n_67, n_626, n_1846);
  xnor g463 (n_70, n_611, n_1837);
  nand g502 (n_661, n_647, n_1790);
  nor g503 (n_652, n_649, n_650);
  nor g506 (n_664, n_654, n_650);
  nor g507 (n_658, n_655, n_656);
  nor g510 (n_672, n_660, n_656);
  nand g513 (n_685, n_649, n_1864);
  nand g514 (n_666, n_664, n_661);
  nand g515 (n_674, n_1854, n_666);
  nor g516 (n_670, n_667, n_668);
  nand g523 (n_689, n_655, n_1882);
  nand g524 (n_677, n_672, n_674);
  nand g525 (n_691, n_668, n_677);
  nand g528 (n_643, n_1878, n_1879);
  xnor g530 (n_83, n_645, n_1791);
  xnor g532 (n_85, n_661, n_1861);
  xnor g535 (n_88, n_685, n_1865);
  xnor g537 (n_91, n_674, n_1870);
  xnor g540 (n_94, n_689, n_1873);
  xnor g542 (n_97, n_691, n_1858);
  nand g569 (n_723, n_706, n_703);
  nor g570 (n_711, n_708, n_709);
  nor g573 (n_726, n_713, n_709);
  nor g574 (n_717, n_714, n_715);
  nor g577 (n_732, n_719, n_715);
  nor g578 (n_721, n_720, B[6]);
  nor g579 (n_734, n_722, B[6]);
  nand g582 (n_752, n_708, n_1866);
  nand g583 (n_728, n_726, n_723);
  nand g584 (n_737, n_1856, n_728);
  nor g592 (n_747, n_1876, n_721);
  nand g593 (n_745, n_732, n_734);
  nand g596 (n_756, n_714, n_1883);
  nand g597 (n_740, n_732, n_737);
  nand g598 (n_758, n_729, n_740);
  nand g604 (n_702, n_747, n_1880);
  xnor g608 (n_86, n_723, n_1862);
  xnor g611 (n_89, n_752, n_1867);
  xnor g613 (n_92, n_737, n_1871);
  xnor g616 (n_95, n_756, n_1874);
  xnor g618 (n_98, n_758, n_1859);
  nand g645 (n_790, n_773, n_1811);
  nor g646 (n_778, n_775, n_776);
  nor g649 (n_793, n_780, n_776);
  nor g650 (n_784, n_781, n_782);
  nor g653 (n_799, n_786, n_782);
  nor g654 (n_788, n_787, n_40);
  nor g655 (n_801, n_789, n_40);
  nand g658 (n_821, n_775, n_1868);
  nand g659 (n_795, n_793, n_790);
  nand g660 (n_804, n_1857, n_795);
  nor g668 (n_814, n_1877, n_788);
  nand g669 (n_812, n_799, n_801);
  nand g672 (n_825, n_781, n_1884);
  nand g673 (n_807, n_799, n_804);
  nand g674 (n_827, n_796, n_807);
  nand g680 (n_816, n_814, n_1881);
  xnor g684 (n_84, n_645, n_1812);
  xnor g686 (n_87, n_790, n_1863);
  xnor g689 (n_90, n_821, n_1869);
  xnor g691 (n_93, n_804, n_1872);
  xnor g694 (n_96, n_825, n_1875);
  xnor g696 (n_99, n_827, n_1860);
  nand g732 (n_859, n_843, n_1793);
  nor g733 (n_848, n_845, n_846);
  nor g736 (n_862, n_850, n_846);
  nor g737 (n_854, n_851, n_852);
  nor g740 (n_868, n_856, n_852);
  nand g744 (n_887, n_845, n_1902);
  nand g745 (n_864, n_862, n_859);
  nand g746 (n_873, n_1890, n_864);
  nor g751 (n_871, n_865, n_858);
  nand g757 (n_891, n_851, n_1922);
  nand g758 (n_876, n_868, n_873);
  nand g759 (n_893, n_865, n_876);
  nand g763 (n_882, n_1916, n_1917);
  xnor g766 (n_120, n_841, n_1794);
  xnor g768 (n_123, n_859, n_1899);
  xnor g771 (n_126, n_887, n_1903);
  xnor g773 (n_129, n_873, n_1908);
  xnor g776 (n_132, n_891, n_1911);
  xnor g778 (n_135, n_893, n_1896);
  nand g812 (n_931, n_911, n_908);
  nor g813 (n_916, n_913, n_914);
  nor g816 (n_934, n_918, n_914);
  nor g817 (n_922, n_919, n_920);
  nor g820 (n_940, n_924, n_920);
  nor g821 (n_928, n_925, n_926);
  nor g824 (n_942, n_930, n_926);
  nand g827 (n_964, n_913, n_1904);
  nand g828 (n_936, n_934, n_931);
  nand g829 (n_947, n_1893, n_936);
  nand g839 (n_955, n_940, n_942);
  nand g842 (n_968, n_919, n_1923);
  nand g843 (n_950, n_940, n_947);
  nand g844 (n_970, n_937, n_950);
  nand g850 (n_959, n_1918, n_1919);
  xnor g855 (n_124, n_931, n_1900);
  xnor g858 (n_127, n_964, n_1905);
  xnor g860 (n_130, n_947, n_1909);
  xnor g863 (n_133, n_968, n_1912);
  xnor g865 (n_136, n_970, n_1897);
  nand g904 (n_1011, n_991, n_1813);
  nor g905 (n_996, n_993, n_994);
  nor g908 (n_1014, n_998, n_994);
  nor g909 (n_1002, n_999, n_1000);
  nor g912 (n_1020, n_1004, n_1000);
  nor g913 (n_1008, n_1005, n_1006);
  nor g916 (n_1022, n_1010, n_1006);
  nand g919 (n_1047, n_993, n_1906);
  nand g920 (n_1016, n_1014, n_1011);
  nand g921 (n_1027, n_1895, n_1016);
  nand g931 (n_1035, n_1020, n_1022);
  nand g934 (n_1051, n_999, n_1924);
  nand g935 (n_1030, n_1020, n_1027);
  nand g936 (n_1053, n_1017, n_1030);
  nand g942 (n_1040, n_1920, n_1921);
  nand g945 (n_151, n_1886, n_1925);
  xnor g947 (n_122, n_841, n_1814);
  xnor g949 (n_125, n_1011, n_1901);
  xnor g952 (n_128, n_1047, n_1907);
  xnor g954 (n_131, n_1027, n_1910);
  xnor g957 (n_134, n_1051, n_1913);
  xnor g959 (n_137, n_1053, n_1898);
  nand g1000 (n_1088, n_1072, n_1796);
  nor g1001 (n_1077, n_1074, n_1075);
  nor g1004 (n_1091, n_1079, n_1075);
  nor g1005 (n_1083, n_1080, n_1081);
  nor g1008 (n_1097, n_1085, n_1081);
  nand g1012 (n_1116, n_1074, n_1943);
  nand g1013 (n_1093, n_1091, n_1088);
  nand g1014 (n_1102, n_1931, n_1093);
  nor g1019 (n_1100, n_1094, n_1087);
  nand g1025 (n_1120, n_1080, n_1963);
  nand g1026 (n_1105, n_1097, n_1102);
  nand g1027 (n_1122, n_1094, n_1105);
  nand g1031 (n_1111, n_1957, n_1958);
  xnor g1034 (n_165, n_1070, n_1797);
  xnor g1036 (n_168, n_1088, n_1940);
  xnor g1039 (n_171, n_1116, n_1944);
  xnor g1041 (n_174, n_1102, n_1949);
  xnor g1044 (n_177, n_1120, n_1952);
  xnor g1046 (n_180, n_1122, n_1937);
  nand g1080 (n_1160, n_1140, n_1137);
  nor g1081 (n_1145, n_1142, n_1143);
  nor g1084 (n_1163, n_1147, n_1143);
  nor g1085 (n_1151, n_1148, n_1149);
  nor g1088 (n_1169, n_1153, n_1149);
  nor g1089 (n_1157, n_1154, n_1155);
  nor g1092 (n_1171, n_1159, n_1155);
  nand g1095 (n_1193, n_1142, n_1945);
  nand g1096 (n_1165, n_1163, n_1160);
  nand g1097 (n_1176, n_1934, n_1165);
  nand g1107 (n_1184, n_1169, n_1171);
  nand g1110 (n_1197, n_1148, n_1964);
  nand g1111 (n_1179, n_1169, n_1176);
  nand g1112 (n_1199, n_1166, n_1179);
  nand g1118 (n_1188, n_1959, n_1960);
  xnor g1123 (n_169, n_1160, n_1941);
  xnor g1126 (n_172, n_1193, n_1946);
  xnor g1128 (n_175, n_1176, n_1950);
  xnor g1131 (n_178, n_1197, n_1953);
  xnor g1133 (n_181, n_1199, n_1938);
  nand g1172 (n_1240, n_1220, n_1815);
  nor g1173 (n_1225, n_1222, n_1223);
  nor g1176 (n_1243, n_1227, n_1223);
  nor g1177 (n_1231, n_1228, n_1229);
  nor g1180 (n_1249, n_1233, n_1229);
  nor g1181 (n_1237, n_1234, n_1235);
  nor g1184 (n_1251, n_1239, n_1235);
  nand g1187 (n_1276, n_1222, n_1947);
  nand g1188 (n_1245, n_1243, n_1240);
  nand g1189 (n_1256, n_1936, n_1245);
  nand g1199 (n_1264, n_1249, n_1251);
  nand g1202 (n_1280, n_1228, n_1965);
  nand g1203 (n_1259, n_1249, n_1256);
  nand g1204 (n_1282, n_1246, n_1259);
  nand g1210 (n_1269, n_1961, n_1962);
  nand g1213 (n_196, n_1927, n_1966);
  xnor g1215 (n_167, n_1070, n_1816);
  xnor g1217 (n_170, n_1240, n_1942);
  xnor g1220 (n_173, n_1276, n_1948);
  xnor g1222 (n_176, n_1256, n_1951);
  xnor g1225 (n_179, n_1280, n_1954);
  xnor g1227 (n_182, n_1282, n_1939);
  nand g1268 (n_1317, n_1301, n_1799);
  nor g1269 (n_1306, n_1303, n_1304);
  nor g1272 (n_1320, n_1308, n_1304);
  nor g1273 (n_1312, n_1309, n_1310);
  nor g1276 (n_1326, n_1314, n_1310);
  nand g1280 (n_1345, n_1303, n_1984);
  nand g1281 (n_1322, n_1320, n_1317);
  nand g1282 (n_1331, n_1972, n_1322);
  nor g1287 (n_1329, n_1323, n_1316);
  nand g1293 (n_1349, n_1309, n_2004);
  nand g1294 (n_1334, n_1326, n_1331);
  nand g1295 (n_1351, n_1323, n_1334);
  nand g1299 (n_1340, n_1998, n_1999);
  xnor g1302 (n_210, n_1299, n_1800);
  xnor g1304 (n_213, n_1317, n_1981);
  xnor g1307 (n_216, n_1345, n_1985);
  xnor g1309 (n_219, n_1331, n_1990);
  xnor g1312 (n_222, n_1349, n_1993);
  xnor g1314 (n_225, n_1351, n_1978);
  nand g1348 (n_1389, n_1369, n_1366);
  nor g1349 (n_1374, n_1371, n_1372);
  nor g1352 (n_1392, n_1376, n_1372);
  nor g1353 (n_1380, n_1377, n_1378);
  nor g1356 (n_1398, n_1382, n_1378);
  nor g1357 (n_1386, n_1383, n_1384);
  nor g1360 (n_1400, n_1388, n_1384);
  nand g1363 (n_1422, n_1371, n_1986);
  nand g1364 (n_1394, n_1392, n_1389);
  nand g1365 (n_1405, n_1975, n_1394);
  nand g1375 (n_1413, n_1398, n_1400);
  nand g1378 (n_1426, n_1377, n_2005);
  nand g1379 (n_1408, n_1398, n_1405);
  nand g1380 (n_1428, n_1395, n_1408);
  nand g1386 (n_1417, n_2000, n_2001);
  xnor g1391 (n_214, n_1389, n_1982);
  xnor g1394 (n_217, n_1422, n_1987);
  xnor g1396 (n_220, n_1405, n_1991);
  xnor g1399 (n_223, n_1426, n_1994);
  xnor g1401 (n_226, n_1428, n_1979);
  nand g1440 (n_1469, n_1449, n_1817);
  nor g1441 (n_1454, n_1451, n_1452);
  nor g1444 (n_1472, n_1456, n_1452);
  nor g1445 (n_1460, n_1457, n_1458);
  nor g1448 (n_1478, n_1462, n_1458);
  nor g1449 (n_1466, n_1463, n_1464);
  nor g1452 (n_1480, n_1468, n_1464);
  nand g1455 (n_1505, n_1451, n_1988);
  nand g1456 (n_1474, n_1472, n_1469);
  nand g1457 (n_1485, n_1977, n_1474);
  nand g1467 (n_1493, n_1478, n_1480);
  nand g1470 (n_1509, n_1457, n_2006);
  nand g1471 (n_1488, n_1478, n_1485);
  nand g1472 (n_1511, n_1475, n_1488);
  nand g1478 (n_1498, n_2002, n_2003);
  nand g1481 (n_241, n_1968, n_2007);
  xnor g1483 (n_212, n_1299, n_1818);
  xnor g1485 (n_215, n_1469, n_1983);
  xnor g1488 (n_218, n_1505, n_1989);
  xnor g1490 (n_221, n_1485, n_1992);
  xnor g1493 (n_224, n_1509, n_1995);
  xnor g1495 (n_227, n_1511, n_1980);
  nand g1536 (n_1546, n_1530, n_1802);
  nor g1537 (n_1535, n_1532, n_1533);
  nor g1540 (n_1549, n_1537, n_1533);
  nor g1541 (n_1541, n_1538, n_1539);
  nor g1544 (n_1555, n_1543, n_1539);
  nand g1548 (n_1574, n_1532, n_2019);
  nand g1549 (n_1551, n_1549, n_1546);
  nand g1550 (n_1560, n_2013, n_1551);
  nor g1555 (n_1558, n_1552, n_1545);
  nand g1561 (n_1578, n_1538, n_2045);
  nand g1562 (n_1563, n_1555, n_1560);
  nand g1563 (n_1580, n_1552, n_1563);
  nand g1567 (n_1569, n_2039, n_2040);
  xnor g1570 (n_255, n_1528, n_1803);
  xnor g1572 (n_258, n_1546, n_2020);
  xnor g1575 (n_261, n_1574, n_2021);
  xnor g1577 (n_264, n_1560, n_2022);
  xnor g1580 (n_267, n_1578, n_2023);
  xnor g1582 (n_270, n_1580, n_2024);
  nand g1616 (n_1618, n_1598, n_1595);
  nor g1617 (n_1603, n_1600, n_1601);
  nor g1620 (n_1621, n_1605, n_1601);
  nor g1621 (n_1609, n_1606, n_1607);
  nor g1624 (n_1627, n_1611, n_1607);
  nor g1625 (n_1615, n_1612, n_1613);
  nor g1628 (n_1629, n_1617, n_1613);
  nand g1631 (n_1651, n_1600, n_2025);
  nand g1632 (n_1623, n_1621, n_1618);
  nand g1633 (n_1634, n_2016, n_1623);
  nand g1643 (n_1642, n_1627, n_1629);
  nand g1646 (n_1655, n_1606, n_2046);
  nand g1647 (n_1637, n_1627, n_1634);
  nand g1648 (n_1657, n_1624, n_1637);
  nand g1654 (n_1646, n_2041, n_2042);
  xnor g1659 (n_259, n_1618, n_2026);
  xnor g1662 (n_262, n_1651, n_2027);
  xnor g1664 (n_265, n_1634, n_2028);
  xnor g1667 (n_268, n_1655, n_2029);
  xnor g1669 (n_271, n_1657, n_2030);
  nand g1708 (n_1698, n_1678, n_1819);
  nor g1709 (n_1683, n_1680, n_1681);
  nor g1712 (n_1701, n_1685, n_1681);
  nor g1713 (n_1689, n_1686, n_1687);
  nor g1716 (n_1707, n_1691, n_1687);
  nor g1717 (n_1695, n_1692, n_1693);
  nor g1720 (n_1709, n_1697, n_1693);
  nand g1723 (n_1734, n_1680, n_2031);
  nand g1724 (n_1703, n_1701, n_1698);
  nand g1725 (n_1714, n_2018, n_1703);
  nand g1735 (n_1722, n_1707, n_1709);
  nand g1738 (n_1738, n_1686, n_2047);
  nand g1739 (n_1717, n_1707, n_1714);
  nand g1740 (n_1740, n_1704, n_1717);
  nand g1746 (n_1727, n_2043, n_2044);
  nand g1749 (n_286, n_2009, n_2048);
  xnor g1751 (n_257, n_1528, n_1820);
  xnor g1753 (n_260, n_1698, n_2032);
  xnor g1756 (n_263, n_1734, n_2033);
  xnor g1758 (n_266, n_1714, n_2034);
  xnor g1761 (n_269, n_1738, n_2035);
  xnor g1763 (n_272, n_1740, n_2036);
  or g1781 (n_1750, wc, A[14]);
  not gc (wc, B[0]);
  or g1782 (n_1751, B[6], wc0);
  not gc0 (wc0, n_353);
  xnor g1783 (n_1752, A[14], B[0]);
  or g1784 (n_372, B[1], wc1);
  not gc1 (wc1, A[13]);
  or g1785 (n_370, wc2, A[12]);
  not gc2 (wc2, B[0]);
  and g1786 (n_1753, B[1], wc3);
  not gc3 (wc3, A[13]);
  or g1787 (n_404, B[0], wc4);
  not gc4 (wc4, A[13]);
  and g1788 (n_401, B[0], wc5);
  not gc5 (wc5, A[13]);
  xnor g1789 (n_1754, A[12], B[0]);
  or g1790 (n_484, B[1], wc6);
  not gc6 (wc6, A[11]);
  or g1791 (n_482, wc7, A[10]);
  not gc7 (wc7, B[0]);
  and g1792 (n_1755, B[1], wc8);
  not gc8 (wc8, A[11]);
  or g1793 (n_532, B[0], wc9);
  not gc9 (wc9, A[11]);
  and g1794 (n_529, B[0], wc10);
  not gc10 (wc10, A[11]);
  xnor g1795 (n_1756, A[10], B[0]);
  or g1796 (n_647, B[1], wc11);
  not gc11 (wc11, A[9]);
  or g1797 (n_645, wc12, A[8]);
  not gc12 (wc12, B[0]);
  and g1798 (n_1757, B[1], wc13);
  not gc13 (wc13, A[9]);
  or g1799 (n_706, B[0], wc14);
  not gc14 (wc14, A[9]);
  and g1800 (n_703, B[0], wc15);
  not gc15 (wc15, A[9]);
  xnor g1801 (n_1758, A[8], B[0]);
  or g1802 (n_843, B[1], wc16);
  not gc16 (wc16, A[7]);
  or g1803 (n_841, wc17, A[6]);
  not gc17 (wc17, B[0]);
  and g1804 (n_1759, B[1], wc18);
  not gc18 (wc18, A[7]);
  or g1805 (n_911, B[0], wc19);
  not gc19 (wc19, A[7]);
  and g1806 (n_908, B[0], wc20);
  not gc20 (wc20, A[7]);
  xnor g1807 (n_1760, A[6], B[0]);
  or g1808 (n_1072, B[1], wc21);
  not gc21 (wc21, A[5]);
  or g1809 (n_1070, wc22, A[4]);
  not gc22 (wc22, B[0]);
  and g1810 (n_1761, B[1], wc23);
  not gc23 (wc23, A[5]);
  or g1811 (n_1140, B[0], wc24);
  not gc24 (wc24, A[5]);
  and g1812 (n_1137, B[0], wc25);
  not gc25 (wc25, A[5]);
  xnor g1813 (n_1762, A[4], B[0]);
  or g1814 (n_1301, B[1], wc26);
  not gc26 (wc26, A[3]);
  or g1815 (n_1299, wc27, A[2]);
  not gc27 (wc27, B[0]);
  and g1816 (n_1763, B[1], wc28);
  not gc28 (wc28, A[3]);
  or g1817 (n_1369, B[0], wc29);
  not gc29 (wc29, A[3]);
  and g1818 (n_1366, B[0], wc30);
  not gc30 (wc30, A[3]);
  xnor g1819 (n_1764, A[2], B[0]);
  or g1820 (n_1530, B[1], wc31);
  not gc31 (wc31, A[1]);
  or g1821 (n_1528, wc32, A[0]);
  not gc32 (wc32, B[0]);
  and g1822 (n_1765, B[1], wc33);
  not gc33 (wc33, A[1]);
  or g1823 (n_1598, B[0], wc34);
  not gc34 (wc34, A[1]);
  and g1824 (n_1595, B[0], wc35);
  not gc35 (wc35, A[1]);
  xnor g1825 (n_1766, A[0], B[0]);
  or g1826 (n_1767, B[1], wc36);
  not gc36 (wc36, n_1750);
  or g1827 (n_1768, wc37, n_298);
  not gc37 (wc37, n_301);
  or g1828 (n_1769, n_295, n_298);
  or g1829 (n_1770, n_351, wc38);
  not gc38 (wc38, n_303);
  or g1830 (n_441, wc39, n_342);
  not gc39 (wc39, A[13]);
  and g1831 (n_1771, wc40, n_342);
  not gc40 (wc40, A[13]);
  or g1832 (n_1772, n_304, wc41);
  not gc41 (wc41, n_305);
  and g1833 (n_1773, wc42, n_305);
  not gc42 (wc42, n_306);
  or g1834 (n_1774, n_353, wc43);
  not gc43 (wc43, n_309);
  or g1835 (n_1775, n_310, wc44);
  not gc44 (wc44, n_311);
  and g1836 (n_322, wc45, n_311);
  not gc45 (wc45, n_312);
  or g1837 (n_587, wc46, n_342);
  not gc46 (wc46, A[11]);
  and g1838 (n_1776, wc47, n_342);
  not gc47 (wc47, A[11]);
  or g1839 (n_773, wc48, n_342);
  not gc48 (wc48, A[9]);
  and g1840 (n_1777, wc49, n_342);
  not gc49 (wc49, A[9]);
  or g1841 (n_991, wc50, n_342);
  not gc50 (wc50, A[7]);
  and g1842 (n_1778, wc51, n_342);
  not gc51 (wc51, A[7]);
  or g1843 (n_1220, wc52, n_342);
  not gc52 (wc52, A[5]);
  and g1844 (n_1779, wc53, n_342);
  not gc53 (wc53, A[5]);
  or g1845 (n_1449, wc54, n_342);
  not gc54 (wc54, A[3]);
  and g1846 (n_1780, wc55, n_342);
  not gc55 (wc55, A[3]);
  or g1847 (n_1678, wc56, n_342);
  not gc56 (wc56, A[1]);
  and g1848 (n_1781, wc57, n_342);
  not gc57 (wc57, A[1]);
  or g1849 (n_1782, n_1753, wc58);
  not gc58 (wc58, n_370);
  xor g1850 (n_1783, n_295, n_1768);
  and g1851 (n_1784, B[6], wc59);
  not gc59 (wc59, n_322);
  or g1852 (n_1785, n_1753, wc60);
  not gc60 (wc60, n_372);
  or g1853 (n_1786, n_401, wc61);
  not gc61 (wc61, n_404);
  or g1854 (n_1787, n_1755, wc62);
  not gc62 (wc62, n_482);
  or g1855 (n_1788, n_1755, wc63);
  not gc63 (wc63, n_484);
  or g1856 (n_1789, n_529, wc64);
  not gc64 (wc64, n_532);
  or g1857 (n_1790, n_1757, wc65);
  not gc65 (wc65, n_645);
  or g1858 (n_1791, n_1757, wc66);
  not gc66 (wc66, n_647);
  or g1859 (n_1792, n_703, wc67);
  not gc67 (wc67, n_706);
  or g1860 (n_1793, n_1759, wc68);
  not gc68 (wc68, n_841);
  or g1861 (n_1794, n_1759, wc69);
  not gc69 (wc69, n_843);
  or g1862 (n_1795, n_908, wc70);
  not gc70 (wc70, n_911);
  or g1863 (n_1796, n_1761, wc71);
  not gc71 (wc71, n_1070);
  or g1864 (n_1797, n_1761, wc72);
  not gc72 (wc72, n_1072);
  or g1865 (n_1798, n_1137, wc73);
  not gc73 (wc73, n_1140);
  or g1866 (n_1799, n_1763, wc74);
  not gc74 (wc74, n_1299);
  or g1867 (n_1800, n_1763, wc75);
  not gc75 (wc75, n_1301);
  or g1868 (n_1801, n_1366, wc76);
  not gc76 (wc76, n_1369);
  or g1869 (n_1802, n_1765, wc77);
  not gc77 (wc77, n_1528);
  or g1870 (n_1803, n_1765, wc78);
  not gc78 (wc78, n_1530);
  or g1871 (n_1804, n_1595, wc79);
  not gc79 (wc79, n_1598);
  or g1872 (n_1805, n_1767, wc80);
  not gc80 (wc80, n_351);
  or g1873 (n_1806, n_1771, wc81);
  not gc81 (wc81, n_370);
  or g1874 (n_1807, n_351, wc82);
  not gc82 (wc82, n_315);
  or g1875 (n_1808, n_1771, wc83);
  not gc83 (wc83, n_441);
  or g1876 (n_1809, n_1776, wc84);
  not gc84 (wc84, n_482);
  or g1877 (n_1810, n_1776, wc85);
  not gc85 (wc85, n_587);
  or g1878 (n_1811, n_1777, wc86);
  not gc86 (wc86, n_645);
  or g1879 (n_1812, n_1777, wc87);
  not gc87 (wc87, n_773);
  or g1880 (n_1813, n_1778, wc88);
  not gc88 (wc88, n_841);
  or g1881 (n_1814, n_1778, wc89);
  not gc89 (wc89, n_991);
  or g1882 (n_1815, n_1779, wc90);
  not gc90 (wc90, n_1070);
  or g1883 (n_1816, n_1779, wc91);
  not gc91 (wc91, n_1220);
  or g1884 (n_1817, n_1780, wc92);
  not gc92 (wc92, n_1299);
  or g1885 (n_1818, n_1780, wc93);
  not gc93 (wc93, n_1449);
  or g1886 (n_1819, n_1781, wc94);
  not gc94 (wc94, n_1528);
  or g1887 (n_1820, n_1781, wc95);
  not gc95 (wc95, n_1678);
  or g1888 (n_32, n_1751, n_1805);
  or g1889 (n_1821, n_353, wc96);
  not gc96 (wc96, n_325);
  or g1890 (n_1822, n_329, wc97);
  not gc97 (wc97, n_325);
  or g1891 (n_1823, wc98, n_1784);
  not gc98 (wc98, n_1822);
  or g1892 (n_34, wc99, wc102);
  and gc102 (wc102, A[14], n_32);
  and gc101 (wc99, wc100, wc101);
  not gc100 (wc101, n_1752);
  not gc99 (wc100, n_32);
  xor g1893 (n_40, n_341, B[6]);
  or g1894 (n_374, B[2], wc103);
  not gc103 (wc103, n_34);
  and g1895 (n_376, B[2], wc104);
  not gc104 (wc104, n_34);
  or g1896 (n_406, B[1], wc105);
  not gc105 (wc105, n_34);
  and g1897 (n_408, B[1], wc106);
  not gc106 (wc106, n_34);
  or g1898 (n_443, wc107, n_1783);
  not gc107 (wc107, n_34);
  and g1899 (n_445, wc108, n_1783);
  not gc108 (wc108, n_34);
  or g1900 (n_1824, n_376, wc109);
  not gc109 (wc109, n_374);
  or g1901 (n_1825, n_408, wc110);
  not gc110 (wc110, n_406);
  or g1902 (n_1826, n_445, wc111);
  not gc111 (wc111, n_443);
  or g1903 (n_1827, wc112, n_375);
  not gc112 (wc112, n_381);
  or g1904 (n_1828, wc113, n_407);
  not gc113 (wc113, n_413);
  or g1905 (n_1829, wc114, n_444);
  not gc114 (wc114, n_450);
  or g1906 (n_48, wc115, n_1751);
  not gc115 (wc115, n_1827);
  or g1907 (n_50, wc116, n_424);
  not gc116 (wc116, n_1828);
  or g1908 (n_1830, wc117, n_461);
  not gc117 (wc117, n_1829);
  and g1909 (n_51, n_50, wc118);
  not gc118 (wc118, n_48);
  or g1910 (n_53, n_1823, n_1830);
  and g1911 (n_54, n_53, wc119);
  not gc119 (wc119, n_50);
  or g1912 (n_58, wc120, wc121, wc122, wc123);
  and gc124 (wc123, wc124, n_47);
  not gc123 (wc124, n_53);
  and gc122 (wc122, n_54, n_46);
  and gc121 (wc121, n_51, n_45);
  and gc120 (wc120, n_48, n_34);
  or g1913 (n_56, wc125, wc126, wc128, wc129);
  and gc131 (wc129, wc130, wc131);
  not gc130 (wc131, n_1754);
  not gc129 (wc130, n_53);
  and gc128 (wc128, A[12], n_54);
  and gc127 (wc126, n_51, wc127);
  not gc126 (wc127, n_1754);
  and gc125 (wc125, A[12], n_48);
  or g1914 (n_57, wc132, wc133, wc134, wc135);
  and gc136 (wc135, wc136, n_44);
  not gc135 (wc136, n_53);
  and gc134 (wc134, n_54, n_1786);
  and gc133 (wc133, n_51, n_43);
  and gc132 (wc132, A[13], n_48);
  or g1915 (n_492, B[4], wc137);
  not gc137 (wc137, n_58);
  or g1916 (n_486, B[2], wc138);
  not gc138 (wc138, n_56);
  and g1917 (n_487, B[3], wc139);
  not gc139 (wc139, n_57);
  or g1918 (n_488, B[3], wc140);
  not gc140 (wc140, n_57);
  and g1919 (n_491, B[2], wc141);
  not gc141 (wc141, n_56);
  and g1920 (n_494, B[4], wc142);
  not gc142 (wc142, n_58);
  or g1921 (n_540, B[3], wc143);
  not gc143 (wc143, n_58);
  or g1922 (n_534, B[1], wc144);
  not gc144 (wc144, n_56);
  and g1923 (n_535, B[2], wc145);
  not gc145 (wc145, n_57);
  or g1924 (n_536, B[2], wc146);
  not gc146 (wc146, n_57);
  and g1925 (n_539, B[1], wc147);
  not gc147 (wc147, n_56);
  and g1926 (n_542, B[3], wc148);
  not gc148 (wc148, n_58);
  or g1927 (n_595, wc149, n_37);
  not gc149 (wc149, n_58);
  or g1928 (n_589, wc150, n_1783);
  not gc150 (wc150, n_56);
  and g1929 (n_590, wc151, n_36);
  not gc151 (wc151, n_57);
  or g1930 (n_591, wc152, n_36);
  not gc152 (wc152, n_57);
  and g1931 (n_594, wc153, n_1783);
  not gc153 (wc153, n_56);
  and g1932 (n_597, wc154, n_37);
  not gc154 (wc154, n_58);
  and g1933 (n_1831, n_488, wc155);
  not gc155 (wc155, n_489);
  or g1934 (n_1832, B[6], wc156);
  not gc156 (wc156, n_503);
  and g1935 (n_1833, n_536, wc157);
  not gc157 (wc157, n_537);
  and g1936 (n_1834, n_591, wc158);
  not gc158 (wc158, n_592);
  or g1937 (n_1835, n_494, wc159);
  not gc159 (wc159, n_492);
  or g1938 (n_1836, n_542, wc160);
  not gc160 (wc160, n_540);
  or g1939 (n_1837, n_597, wc161);
  not gc161 (wc161, n_595);
  or g1940 (n_1838, n_491, wc162);
  not gc162 (wc162, n_486);
  or g1941 (n_1839, n_539, wc163);
  not gc163 (wc163, n_534);
  or g1942 (n_1840, n_594, wc164);
  not gc164 (wc164, n_589);
  or g1943 (n_1841, n_491, wc165);
  not gc165 (wc165, n_495);
  or g1944 (n_1842, wc166, n_487);
  not gc166 (wc166, n_488);
  or g1945 (n_1843, n_539, wc167);
  not gc167 (wc167, n_543);
  or g1946 (n_1844, wc168, n_535);
  not gc168 (wc168, n_536);
  or g1947 (n_1845, n_594, wc169);
  not gc169 (wc169, n_598);
  or g1948 (n_1846, wc170, n_590);
  not gc170 (wc170, n_591);
  and g1949 (n_1847, wc171, n_493);
  not gc171 (wc171, B[6]);
  and g1950 (n_1848, n_310, n_541);
  and g1951 (n_1849, n_453, n_596);
  or g1952 (n_1850, n_1832, wc172);
  not gc172 (wc172, n_505);
  or g1953 (n_1851, n_563, wc173);
  not gc173 (wc173, n_556);
  or g1954 (n_1852, n_618, wc174);
  not gc174 (wc174, n_611);
  or g1955 (n_480, wc175, n_1847);
  not gc175 (wc175, n_1850);
  or g1956 (n_528, wc176, n_1848);
  not gc176 (wc176, n_1851);
  or g1957 (n_1853, wc177, n_1849);
  not gc177 (wc177, n_1852);
  or g1958 (n_74, wc178, n_1823);
  not gc178 (wc178, n_1853);
  and g1959 (n_73, wc179, n_480);
  not gc179 (wc179, n_528);
  or g1960 (n_81, wc180, wc182, wc183, wc184);
  and gc185 (wc184, wc185, n_70);
  not gc184 (wc185, n_74);
  and gc183 (wc183, n_69, n_75);
  and gc182 (wc182, n_73, n_68);
  and gc181 (wc180, wc181, n_58);
  not gc180 (wc181, n_480);
  or g1961 (n_79, wc186, wc188, wc189, wc190);
  and gc191 (wc190, wc191, n_64);
  not gc190 (wc191, n_74);
  and gc189 (wc189, n_63, n_75);
  and gc188 (wc188, n_73, n_62);
  and gc187 (wc186, wc187, n_56);
  not gc186 (wc187, n_480);
  or g1962 (n_80, wc192, wc194, wc195, wc196);
  and gc197 (wc196, wc197, n_67);
  not gc196 (wc197, n_74);
  and gc195 (wc195, n_66, n_75);
  and gc194 (wc194, n_73, n_65);
  and gc193 (wc192, wc193, n_57);
  not gc192 (wc193, n_480);
  or g1963 (n_77, wc198, wc200, wc202, wc203);
  and gc205 (wc203, wc204, wc205);
  not gc204 (wc205, n_1756);
  not gc203 (wc204, n_74);
  and gc202 (wc202, A[10], n_75);
  and gc201 (wc200, n_73, wc201);
  not gc200 (wc201, n_1756);
  and gc199 (wc198, A[10], wc199);
  not gc198 (wc199, n_480);
  or g1964 (n_78, wc206, wc208, wc209, wc210);
  and gc211 (wc210, wc211, n_61);
  not gc210 (wc211, n_74);
  and gc209 (wc209, n_1789, n_75);
  and gc208 (wc208, n_73, n_60);
  and gc207 (wc206, A[11], wc207);
  not gc206 (wc207, n_480);
  and g1965 (n_667, B[6], wc212);
  not gc212 (wc212, n_81);
  or g1966 (n_655, B[4], wc213);
  not gc213 (wc213, n_79);
  and g1967 (n_656, B[5], wc214);
  not gc214 (wc214, n_80);
  or g1968 (n_657, B[5], wc215);
  not gc215 (wc215, n_80);
  or g1969 (n_669, B[6], wc216);
  not gc216 (wc216, n_81);
  or g1970 (n_649, B[2], wc217);
  not gc217 (wc217, n_77);
  and g1971 (n_650, B[3], wc218);
  not gc218 (wc218, n_78);
  or g1972 (n_651, B[3], wc219);
  not gc219 (wc219, n_78);
  and g1973 (n_654, B[2], wc220);
  not gc220 (wc220, n_77);
  and g1974 (n_660, B[4], wc221);
  not gc221 (wc221, n_79);
  or g1975 (n_714, B[3], wc222);
  not gc222 (wc222, n_79);
  and g1976 (n_715, B[4], wc223);
  not gc223 (wc223, n_80);
  or g1977 (n_716, B[4], wc224);
  not gc224 (wc224, n_80);
  and g1978 (n_722, B[5], wc225);
  not gc225 (wc225, n_81);
  or g1979 (n_720, B[5], wc226);
  not gc226 (wc226, n_81);
  or g1980 (n_708, B[1], wc227);
  not gc227 (wc227, n_77);
  and g1981 (n_709, B[2], wc228);
  not gc228 (wc228, n_78);
  or g1982 (n_710, B[2], wc229);
  not gc229 (wc229, n_78);
  and g1983 (n_713, B[1], wc230);
  not gc230 (wc230, n_77);
  and g1984 (n_719, B[3], wc231);
  not gc231 (wc231, n_79);
  or g1985 (n_781, wc232, n_37);
  not gc232 (wc232, n_79);
  and g1986 (n_782, wc233, n_38);
  not gc233 (wc233, n_80);
  or g1987 (n_783, wc234, n_38);
  not gc234 (wc234, n_80);
  and g1988 (n_789, wc235, n_39);
  not gc235 (wc235, n_81);
  or g1989 (n_787, wc236, n_39);
  not gc236 (wc236, n_81);
  or g1990 (n_775, wc237, n_1783);
  not gc237 (wc237, n_77);
  and g1991 (n_776, wc238, n_36);
  not gc238 (wc238, n_78);
  or g1992 (n_777, wc239, n_36);
  not gc239 (wc239, n_78);
  and g1993 (n_780, wc240, n_1783);
  not gc240 (wc240, n_77);
  and g1994 (n_786, wc241, n_37);
  not gc241 (wc241, n_79);
  and g1995 (n_668, n_657, wc242);
  not gc242 (wc242, n_658);
  and g1996 (n_1854, n_651, wc243);
  not gc243 (wc243, n_652);
  or g1997 (n_1855, n_667, wc244);
  not gc244 (wc244, n_672);
  and g1998 (n_729, n_716, wc245);
  not gc245 (wc245, n_717);
  and g1999 (n_1856, n_710, wc246);
  not gc246 (wc246, n_711);
  and g2000 (n_796, n_783, wc247);
  not gc247 (wc247, n_784);
  and g2001 (n_1857, n_777, wc248);
  not gc248 (wc248, n_778);
  or g2002 (n_1858, wc249, n_667);
  not gc249 (wc249, n_669);
  or g2003 (n_1859, wc250, n_722);
  not gc250 (wc250, n_720);
  or g2004 (n_1860, wc251, n_789);
  not gc251 (wc251, n_787);
  or g2005 (n_1861, n_654, wc252);
  not gc252 (wc252, n_649);
  or g2006 (n_1862, n_713, wc253);
  not gc253 (wc253, n_708);
  or g2007 (n_1863, n_780, wc254);
  not gc254 (wc254, n_775);
  or g2008 (n_1864, n_654, wc255);
  not gc255 (wc255, n_661);
  or g2009 (n_1865, wc256, n_650);
  not gc256 (wc256, n_651);
  or g2010 (n_1866, n_713, wc257);
  not gc257 (wc257, n_723);
  or g2011 (n_1867, wc258, n_709);
  not gc258 (wc258, n_710);
  or g2012 (n_1868, n_780, wc259);
  not gc259 (wc259, n_790);
  or g2013 (n_1869, wc260, n_776);
  not gc260 (wc260, n_777);
  or g2014 (n_1870, n_660, wc261);
  not gc261 (wc261, n_655);
  or g2015 (n_1871, n_719, wc262);
  not gc262 (wc262, n_714);
  or g2016 (n_1872, n_786, wc263);
  not gc263 (wc263, n_781);
  or g2017 (n_1873, wc264, n_656);
  not gc264 (wc264, n_657);
  or g2018 (n_1874, wc265, n_715);
  not gc265 (wc265, n_716);
  or g2019 (n_1875, wc266, n_782);
  not gc266 (wc266, n_783);
  and g2020 (n_1876, wc267, n_734);
  not gc267 (wc267, n_729);
  and g2021 (n_1877, wc268, n_801);
  not gc268 (wc268, n_796);
  and g2022 (n_1878, n_669, wc269);
  not gc269 (wc269, n_670);
  or g2023 (n_1879, n_1855, wc270);
  not gc270 (wc270, n_674);
  or g2024 (n_1880, n_745, wc271);
  not gc271 (wc271, n_737);
  or g2025 (n_1881, n_812, wc272);
  not gc272 (wc272, n_804);
  or g2026 (n_1882, n_660, wc273);
  not gc273 (wc273, n_674);
  or g2027 (n_1883, n_719, wc274);
  not gc274 (wc274, n_737);
  or g2028 (n_1884, n_786, wc275);
  not gc275 (wc275, n_804);
  or g2029 (n_104, n_1823, wc276);
  not gc276 (wc276, n_816);
  and g2030 (n_102, wc277, n_643);
  not gc277 (wc277, n_702);
  or g2031 (n_116, wc278, wc280, wc281, wc282);
  and gc283 (wc282, wc283, n_99);
  not gc282 (wc283, n_104);
  and gc281 (wc281, n_98, n_105);
  and gc280 (wc280, n_102, n_97);
  and gc279 (wc278, n_81, wc279);
  not gc278 (wc279, n_643);
  or g2032 (n_112, wc284, wc286, wc287, wc288);
  and gc289 (wc288, wc289, n_87);
  not gc288 (wc289, n_104);
  and gc287 (wc287, n_86, n_105);
  and gc286 (wc286, n_102, n_85);
  and gc285 (wc284, n_77, wc285);
  not gc284 (wc285, n_643);
  or g2033 (n_113, wc290, wc292, wc293, wc294);
  and gc295 (wc294, wc295, n_90);
  not gc294 (wc295, n_104);
  and gc293 (wc293, n_89, n_105);
  and gc292 (wc292, n_102, n_88);
  and gc291 (wc290, n_78, wc291);
  not gc290 (wc291, n_643);
  or g2034 (n_114, wc296, wc298, wc299, wc300);
  and gc301 (wc300, wc301, n_93);
  not gc300 (wc301, n_104);
  and gc299 (wc299, n_92, n_105);
  and gc298 (wc298, n_102, n_91);
  and gc297 (wc296, n_79, wc297);
  not gc296 (wc297, n_643);
  or g2035 (n_115, wc302, wc304, wc305, wc306);
  and gc307 (wc306, wc307, n_96);
  not gc306 (wc307, n_104);
  and gc305 (wc305, n_95, n_105);
  and gc304 (wc304, n_102, n_94);
  and gc303 (wc302, n_80, wc303);
  not gc302 (wc303, n_643);
  or g2036 (n_110, wc308, wc310, wc312, wc313);
  and gc315 (wc313, wc314, wc315);
  not gc314 (wc315, n_1758);
  not gc313 (wc314, n_104);
  and gc312 (wc312, A[8], n_105);
  and gc311 (wc310, n_102, wc311);
  not gc310 (wc311, n_1758);
  and gc309 (wc308, A[8], wc309);
  not gc308 (wc309, n_643);
  or g2037 (n_111, wc316, wc318, wc319, wc320);
  and gc321 (wc320, wc321, n_84);
  not gc320 (wc321, n_104);
  and gc319 (wc319, n_1792, n_105);
  and gc318 (wc318, n_102, n_83);
  and gc317 (wc316, A[9], wc317);
  not gc316 (wc317, n_643);
  or g2038 (n_851, B[4], wc322);
  not gc322 (wc322, n_112);
  and g2039 (n_852, B[5], wc323);
  not gc323 (wc323, n_113);
  or g2040 (n_853, B[5], wc324);
  not gc324 (wc324, n_113);
  and g2041 (n_858, B[6], wc325);
  not gc325 (wc325, n_114);
  or g2042 (n_857, B[6], wc326);
  not gc326 (wc326, n_114);
  or g2043 (n_845, B[2], wc327);
  not gc327 (wc327, n_110);
  and g2044 (n_846, B[3], wc328);
  not gc328 (wc328, n_111);
  or g2045 (n_847, B[3], wc329);
  not gc329 (wc329, n_111);
  and g2046 (n_850, B[2], wc330);
  not gc330 (wc330, n_110);
  and g2047 (n_856, B[4], wc331);
  not gc331 (wc331, n_112);
  or g2048 (n_919, B[3], wc332);
  not gc332 (wc332, n_112);
  and g2049 (n_920, B[4], wc333);
  not gc333 (wc333, n_113);
  or g2050 (n_921, B[4], wc334);
  not gc334 (wc334, n_113);
  and g2051 (n_930, B[5], wc335);
  not gc335 (wc335, n_114);
  and g2052 (n_926, B[6], wc336);
  not gc336 (wc336, n_115);
  or g2053 (n_925, B[5], wc337);
  not gc337 (wc337, n_114);
  or g2054 (n_1885, B[6], wc338);
  not gc338 (wc338, n_115);
  or g2055 (n_913, B[1], wc339);
  not gc339 (wc339, n_110);
  and g2056 (n_914, B[2], wc340);
  not gc340 (wc340, n_111);
  or g2057 (n_915, B[2], wc341);
  not gc341 (wc341, n_111);
  and g2058 (n_918, B[1], wc342);
  not gc342 (wc342, n_110);
  and g2059 (n_924, B[3], wc343);
  not gc343 (wc343, n_112);
  or g2060 (n_1886, wc344, n_1823);
  not gc344 (wc344, n_116);
  or g2061 (n_999, wc345, n_37);
  not gc345 (wc345, n_112);
  and g2062 (n_1000, wc346, n_38);
  not gc346 (wc346, n_113);
  or g2063 (n_1001, wc347, n_38);
  not gc347 (wc347, n_113);
  and g2064 (n_1010, wc348, n_39);
  not gc348 (wc348, n_114);
  and g2065 (n_1006, wc349, n_40);
  not gc349 (wc349, n_115);
  or g2066 (n_1005, wc350, n_39);
  not gc350 (wc350, n_114);
  or g2067 (n_1887, wc351, n_40);
  not gc351 (wc351, n_115);
  or g2068 (n_993, wc352, n_1783);
  not gc352 (wc352, n_110);
  and g2069 (n_994, wc353, n_36);
  not gc353 (wc353, n_111);
  or g2070 (n_995, wc354, n_36);
  not gc354 (wc354, n_111);
  and g2071 (n_998, wc355, n_1783);
  not gc355 (wc355, n_110);
  and g2072 (n_1004, wc356, n_37);
  not gc356 (wc356, n_112);
  and g2073 (n_1888, wc357, n_1823);
  not gc357 (wc357, n_116);
  and g2074 (n_865, n_853, wc358);
  not gc358 (wc358, n_854);
  and g2075 (n_1889, n_857, wc359);
  not gc359 (wc359, n_115);
  and g2076 (n_1890, n_847, wc360);
  not gc360 (wc360, n_848);
  or g2077 (n_1891, n_858, wc361);
  not gc361 (wc361, n_868);
  and g2078 (n_937, n_921, wc362);
  not gc362 (wc362, n_922);
  and g2079 (n_1892, n_1885, wc363);
  not gc363 (wc363, n_928);
  and g2080 (n_1893, n_915, wc364);
  not gc364 (wc364, n_916);
  and g2081 (n_1017, n_1001, wc365);
  not gc365 (wc365, n_1002);
  and g2082 (n_1894, n_1887, wc366);
  not gc366 (wc366, n_1008);
  and g2083 (n_1895, n_995, wc367);
  not gc367 (wc367, n_996);
  or g2084 (n_1896, wc368, n_858);
  not gc368 (wc368, n_857);
  or g2085 (n_1897, wc369, n_930);
  not gc369 (wc369, n_925);
  or g2086 (n_1898, wc370, n_1010);
  not gc370 (wc370, n_1005);
  or g2087 (n_1899, n_850, wc371);
  not gc371 (wc371, n_845);
  or g2088 (n_1900, n_918, wc372);
  not gc372 (wc372, n_913);
  or g2089 (n_1901, n_998, wc373);
  not gc373 (wc373, n_993);
  or g2090 (n_1902, n_850, wc374);
  not gc374 (wc374, n_859);
  or g2091 (n_1903, wc375, n_846);
  not gc375 (wc375, n_847);
  or g2092 (n_1904, n_918, wc376);
  not gc376 (wc376, n_931);
  or g2093 (n_1905, wc377, n_914);
  not gc377 (wc377, n_915);
  or g2094 (n_1906, n_998, wc378);
  not gc378 (wc378, n_1011);
  or g2095 (n_1907, wc379, n_994);
  not gc379 (wc379, n_995);
  or g2096 (n_1908, n_856, wc380);
  not gc380 (wc380, n_851);
  or g2097 (n_1909, n_924, wc381);
  not gc381 (wc381, n_919);
  or g2098 (n_1910, n_1004, wc382);
  not gc382 (wc382, n_999);
  or g2099 (n_1911, wc383, n_852);
  not gc383 (wc383, n_853);
  or g2100 (n_1912, wc384, n_920);
  not gc384 (wc384, n_921);
  or g2101 (n_1913, wc385, n_1000);
  not gc385 (wc385, n_1001);
  and g2102 (n_1914, wc386, n_942);
  not gc386 (wc386, n_937);
  and g2103 (n_1915, wc387, n_1022);
  not gc387 (wc387, n_1017);
  and g2104 (n_1916, n_1889, wc388);
  not gc388 (wc388, n_871);
  or g2105 (n_1917, n_1891, wc389);
  not gc389 (wc389, n_873);
  and g2106 (n_1918, wc390, n_1892);
  not gc390 (wc390, n_1914);
  or g2107 (n_1919, n_955, wc391);
  not gc391 (wc391, n_947);
  and g2108 (n_1920, wc392, n_1894);
  not gc392 (wc392, n_1915);
  or g2109 (n_1921, n_1035, wc393);
  not gc393 (wc393, n_1027);
  or g2110 (n_1922, n_856, wc394);
  not gc394 (wc394, n_873);
  or g2111 (n_1923, n_924, wc395);
  not gc395 (wc395, n_947);
  or g2112 (n_1924, n_1004, wc396);
  not gc396 (wc396, n_1027);
  or g2113 (n_1925, n_1888, wc397);
  not gc397 (wc397, n_1040);
  or g2114 (n_839, n_882, n_116);
  or g2115 (n_907, n_959, n_116);
  and g2116 (n_147, wc398, n_839);
  not gc398 (wc398, n_907);
  and g2117 (n_150, n_907, wc399);
  not gc399 (wc399, n_151);
  or g2118 (n_161, wc400, wc402, wc403, wc404);
  and gc404 (wc404, n_137, n_151);
  and gc403 (wc403, n_150, n_136);
  and gc402 (wc402, n_147, n_135);
  and gc401 (wc400, wc401, n_114);
  not gc400 (wc401, n_839);
  or g2119 (n_157, wc405, wc407, wc408, wc409);
  and gc409 (wc409, n_125, n_151);
  and gc408 (wc408, n_150, n_124);
  and gc407 (wc407, n_147, n_123);
  and gc406 (wc405, wc406, n_110);
  not gc405 (wc406, n_839);
  or g2120 (n_158, wc410, wc412, wc413, wc414);
  and gc414 (wc414, n_128, n_151);
  and gc413 (wc413, n_150, n_127);
  and gc412 (wc412, n_147, n_126);
  and gc411 (wc410, wc411, n_111);
  not gc410 (wc411, n_839);
  or g2121 (n_159, wc415, wc417, wc418, wc419);
  and gc419 (wc419, n_131, n_151);
  and gc418 (wc418, n_150, n_130);
  and gc417 (wc417, n_147, n_129);
  and gc416 (wc415, wc416, n_112);
  not gc415 (wc416, n_839);
  or g2122 (n_160, wc420, wc422, wc423, wc424);
  and gc424 (wc424, n_134, n_151);
  and gc423 (wc423, n_150, n_133);
  and gc422 (wc422, n_147, n_132);
  and gc421 (wc420, wc421, n_113);
  not gc420 (wc421, n_839);
  or g2123 (n_155, wc425, wc427, wc429, wc430);
  and gc431 (wc430, wc431, n_151);
  not gc430 (wc431, n_1760);
  and gc429 (wc429, A[6], n_150);
  and gc428 (wc427, n_147, wc428);
  not gc427 (wc428, n_1760);
  and gc426 (wc425, A[6], wc426);
  not gc425 (wc426, n_839);
  or g2124 (n_156, wc432, wc434, wc435, wc436);
  and gc436 (wc436, n_122, n_151);
  and gc435 (wc435, n_150, n_1795);
  and gc434 (wc434, n_147, n_120);
  and gc433 (wc432, A[7], wc433);
  not gc432 (wc433, n_839);
  or g2125 (n_1080, B[4], wc437);
  not gc437 (wc437, n_157);
  and g2126 (n_1081, B[5], wc438);
  not gc438 (wc438, n_158);
  or g2127 (n_1082, B[5], wc439);
  not gc439 (wc439, n_158);
  and g2128 (n_1087, B[6], wc440);
  not gc440 (wc440, n_159);
  or g2129 (n_1086, B[6], wc441);
  not gc441 (wc441, n_159);
  or g2130 (n_1074, B[2], wc442);
  not gc442 (wc442, n_155);
  and g2131 (n_1075, B[3], wc443);
  not gc443 (wc443, n_156);
  or g2132 (n_1076, B[3], wc444);
  not gc444 (wc444, n_156);
  and g2133 (n_1079, B[2], wc445);
  not gc445 (wc445, n_155);
  and g2134 (n_1085, B[4], wc446);
  not gc446 (wc446, n_157);
  or g2135 (n_1148, B[3], wc447);
  not gc447 (wc447, n_157);
  and g2136 (n_1149, B[4], wc448);
  not gc448 (wc448, n_158);
  or g2137 (n_1150, B[4], wc449);
  not gc449 (wc449, n_158);
  and g2138 (n_1159, B[5], wc450);
  not gc450 (wc450, n_159);
  and g2139 (n_1155, B[6], wc451);
  not gc451 (wc451, n_160);
  or g2140 (n_1154, B[5], wc452);
  not gc452 (wc452, n_159);
  or g2141 (n_1926, B[6], wc453);
  not gc453 (wc453, n_160);
  or g2142 (n_1142, B[1], wc454);
  not gc454 (wc454, n_155);
  and g2143 (n_1143, B[2], wc455);
  not gc455 (wc455, n_156);
  or g2144 (n_1144, B[2], wc456);
  not gc456 (wc456, n_156);
  and g2145 (n_1147, B[1], wc457);
  not gc457 (wc457, n_155);
  and g2146 (n_1153, B[3], wc458);
  not gc458 (wc458, n_157);
  or g2147 (n_1927, wc459, n_1823);
  not gc459 (wc459, n_161);
  or g2148 (n_1228, wc460, n_37);
  not gc460 (wc460, n_157);
  and g2149 (n_1229, wc461, n_38);
  not gc461 (wc461, n_158);
  or g2150 (n_1230, wc462, n_38);
  not gc462 (wc462, n_158);
  and g2151 (n_1239, wc463, n_39);
  not gc463 (wc463, n_159);
  and g2152 (n_1235, wc464, n_40);
  not gc464 (wc464, n_160);
  or g2153 (n_1234, wc465, n_39);
  not gc465 (wc465, n_159);
  or g2154 (n_1928, wc466, n_40);
  not gc466 (wc466, n_160);
  or g2155 (n_1222, wc467, n_1783);
  not gc467 (wc467, n_155);
  and g2156 (n_1223, wc468, n_36);
  not gc468 (wc468, n_156);
  or g2157 (n_1224, wc469, n_36);
  not gc469 (wc469, n_156);
  and g2158 (n_1227, wc470, n_1783);
  not gc470 (wc470, n_155);
  and g2159 (n_1233, wc471, n_37);
  not gc471 (wc471, n_157);
  and g2160 (n_1929, wc472, n_1823);
  not gc472 (wc472, n_161);
  and g2161 (n_1094, n_1082, wc473);
  not gc473 (wc473, n_1083);
  and g2162 (n_1930, n_1086, wc474);
  not gc474 (wc474, n_160);
  and g2163 (n_1931, n_1076, wc475);
  not gc475 (wc475, n_1077);
  or g2164 (n_1932, n_1087, wc476);
  not gc476 (wc476, n_1097);
  and g2165 (n_1166, n_1150, wc477);
  not gc477 (wc477, n_1151);
  and g2166 (n_1933, n_1926, wc478);
  not gc478 (wc478, n_1157);
  and g2167 (n_1934, n_1144, wc479);
  not gc479 (wc479, n_1145);
  and g2168 (n_1246, n_1230, wc480);
  not gc480 (wc480, n_1231);
  and g2169 (n_1935, n_1928, wc481);
  not gc481 (wc481, n_1237);
  and g2170 (n_1936, n_1224, wc482);
  not gc482 (wc482, n_1225);
  or g2171 (n_1937, wc483, n_1087);
  not gc483 (wc483, n_1086);
  or g2172 (n_1938, wc484, n_1159);
  not gc484 (wc484, n_1154);
  or g2173 (n_1939, wc485, n_1239);
  not gc485 (wc485, n_1234);
  or g2174 (n_1940, n_1079, wc486);
  not gc486 (wc486, n_1074);
  or g2175 (n_1941, n_1147, wc487);
  not gc487 (wc487, n_1142);
  or g2176 (n_1942, n_1227, wc488);
  not gc488 (wc488, n_1222);
  or g2177 (n_1943, n_1079, wc489);
  not gc489 (wc489, n_1088);
  or g2178 (n_1944, wc490, n_1075);
  not gc490 (wc490, n_1076);
  or g2179 (n_1945, n_1147, wc491);
  not gc491 (wc491, n_1160);
  or g2180 (n_1946, wc492, n_1143);
  not gc492 (wc492, n_1144);
  or g2181 (n_1947, n_1227, wc493);
  not gc493 (wc493, n_1240);
  or g2182 (n_1948, wc494, n_1223);
  not gc494 (wc494, n_1224);
  or g2183 (n_1949, n_1085, wc495);
  not gc495 (wc495, n_1080);
  or g2184 (n_1950, n_1153, wc496);
  not gc496 (wc496, n_1148);
  or g2185 (n_1951, n_1233, wc497);
  not gc497 (wc497, n_1228);
  or g2186 (n_1952, wc498, n_1081);
  not gc498 (wc498, n_1082);
  or g2187 (n_1953, wc499, n_1149);
  not gc499 (wc499, n_1150);
  or g2188 (n_1954, wc500, n_1229);
  not gc500 (wc500, n_1230);
  and g2189 (n_1955, wc501, n_1171);
  not gc501 (wc501, n_1166);
  and g2190 (n_1956, wc502, n_1251);
  not gc502 (wc502, n_1246);
  and g2191 (n_1957, n_1930, wc503);
  not gc503 (wc503, n_1100);
  or g2192 (n_1958, n_1932, wc504);
  not gc504 (wc504, n_1102);
  and g2193 (n_1959, wc505, n_1933);
  not gc505 (wc505, n_1955);
  or g2194 (n_1960, n_1184, wc506);
  not gc506 (wc506, n_1176);
  and g2195 (n_1961, wc507, n_1935);
  not gc507 (wc507, n_1956);
  or g2196 (n_1962, n_1264, wc508);
  not gc508 (wc508, n_1256);
  or g2197 (n_1963, n_1085, wc509);
  not gc509 (wc509, n_1102);
  or g2198 (n_1964, n_1153, wc510);
  not gc510 (wc510, n_1176);
  or g2199 (n_1965, n_1233, wc511);
  not gc511 (wc511, n_1256);
  or g2200 (n_1966, n_1929, wc512);
  not gc512 (wc512, n_1269);
  or g2201 (n_1068, n_1111, n_161);
  or g2202 (n_1136, n_1188, n_161);
  and g2203 (n_192, wc513, n_1068);
  not gc513 (wc513, n_1136);
  and g2204 (n_195, n_1136, wc514);
  not gc514 (wc514, n_196);
  or g2205 (n_206, wc515, wc517, wc518, wc519);
  and gc519 (wc519, n_182, n_196);
  and gc518 (wc518, n_195, n_181);
  and gc517 (wc517, n_192, n_180);
  and gc516 (wc515, wc516, n_159);
  not gc515 (wc516, n_1068);
  or g2206 (n_202, wc520, wc522, wc523, wc524);
  and gc524 (wc524, n_170, n_196);
  and gc523 (wc523, n_195, n_169);
  and gc522 (wc522, n_192, n_168);
  and gc521 (wc520, wc521, n_155);
  not gc520 (wc521, n_1068);
  or g2207 (n_203, wc525, wc527, wc528, wc529);
  and gc529 (wc529, n_173, n_196);
  and gc528 (wc528, n_195, n_172);
  and gc527 (wc527, n_192, n_171);
  and gc526 (wc525, wc526, n_156);
  not gc525 (wc526, n_1068);
  or g2208 (n_204, wc530, wc532, wc533, wc534);
  and gc534 (wc534, n_176, n_196);
  and gc533 (wc533, n_195, n_175);
  and gc532 (wc532, n_192, n_174);
  and gc531 (wc530, wc531, n_157);
  not gc530 (wc531, n_1068);
  or g2209 (n_205, wc535, wc537, wc538, wc539);
  and gc539 (wc539, n_179, n_196);
  and gc538 (wc538, n_195, n_178);
  and gc537 (wc537, n_192, n_177);
  and gc536 (wc535, wc536, n_158);
  not gc535 (wc536, n_1068);
  or g2210 (n_200, wc540, wc542, wc544, wc545);
  and gc546 (wc545, wc546, n_196);
  not gc545 (wc546, n_1762);
  and gc544 (wc544, A[4], n_195);
  and gc543 (wc542, n_192, wc543);
  not gc542 (wc543, n_1762);
  and gc541 (wc540, A[4], wc541);
  not gc540 (wc541, n_1068);
  or g2211 (n_201, wc547, wc549, wc550, wc551);
  and gc551 (wc551, n_167, n_196);
  and gc550 (wc550, n_195, n_1798);
  and gc549 (wc549, n_192, n_165);
  and gc548 (wc547, A[5], wc548);
  not gc547 (wc548, n_1068);
  or g2212 (n_1309, B[4], wc552);
  not gc552 (wc552, n_202);
  and g2213 (n_1310, B[5], wc553);
  not gc553 (wc553, n_203);
  or g2214 (n_1311, B[5], wc554);
  not gc554 (wc554, n_203);
  and g2215 (n_1316, B[6], wc555);
  not gc555 (wc555, n_204);
  or g2216 (n_1315, B[6], wc556);
  not gc556 (wc556, n_204);
  or g2217 (n_1303, B[2], wc557);
  not gc557 (wc557, n_200);
  and g2218 (n_1304, B[3], wc558);
  not gc558 (wc558, n_201);
  or g2219 (n_1305, B[3], wc559);
  not gc559 (wc559, n_201);
  and g2220 (n_1308, B[2], wc560);
  not gc560 (wc560, n_200);
  and g2221 (n_1314, B[4], wc561);
  not gc561 (wc561, n_202);
  or g2222 (n_1377, B[3], wc562);
  not gc562 (wc562, n_202);
  and g2223 (n_1378, B[4], wc563);
  not gc563 (wc563, n_203);
  or g2224 (n_1379, B[4], wc564);
  not gc564 (wc564, n_203);
  and g2225 (n_1388, B[5], wc565);
  not gc565 (wc565, n_204);
  and g2226 (n_1384, B[6], wc566);
  not gc566 (wc566, n_205);
  or g2227 (n_1383, B[5], wc567);
  not gc567 (wc567, n_204);
  or g2228 (n_1967, B[6], wc568);
  not gc568 (wc568, n_205);
  or g2229 (n_1371, B[1], wc569);
  not gc569 (wc569, n_200);
  and g2230 (n_1372, B[2], wc570);
  not gc570 (wc570, n_201);
  or g2231 (n_1373, B[2], wc571);
  not gc571 (wc571, n_201);
  and g2232 (n_1376, B[1], wc572);
  not gc572 (wc572, n_200);
  and g2233 (n_1382, B[3], wc573);
  not gc573 (wc573, n_202);
  or g2234 (n_1968, wc574, n_1823);
  not gc574 (wc574, n_206);
  or g2235 (n_1457, wc575, n_37);
  not gc575 (wc575, n_202);
  and g2236 (n_1458, wc576, n_38);
  not gc576 (wc576, n_203);
  or g2237 (n_1459, wc577, n_38);
  not gc577 (wc577, n_203);
  and g2238 (n_1468, wc578, n_39);
  not gc578 (wc578, n_204);
  and g2239 (n_1464, wc579, n_40);
  not gc579 (wc579, n_205);
  or g2240 (n_1463, wc580, n_39);
  not gc580 (wc580, n_204);
  or g2241 (n_1969, wc581, n_40);
  not gc581 (wc581, n_205);
  or g2242 (n_1451, wc582, n_1783);
  not gc582 (wc582, n_200);
  and g2243 (n_1452, wc583, n_36);
  not gc583 (wc583, n_201);
  or g2244 (n_1453, wc584, n_36);
  not gc584 (wc584, n_201);
  and g2245 (n_1456, wc585, n_1783);
  not gc585 (wc585, n_200);
  and g2246 (n_1462, wc586, n_37);
  not gc586 (wc586, n_202);
  and g2247 (n_1970, wc587, n_1823);
  not gc587 (wc587, n_206);
  and g2248 (n_1323, n_1311, wc588);
  not gc588 (wc588, n_1312);
  and g2249 (n_1971, n_1315, wc589);
  not gc589 (wc589, n_205);
  and g2250 (n_1972, n_1305, wc590);
  not gc590 (wc590, n_1306);
  or g2251 (n_1973, n_1316, wc591);
  not gc591 (wc591, n_1326);
  and g2252 (n_1395, n_1379, wc592);
  not gc592 (wc592, n_1380);
  and g2253 (n_1974, n_1967, wc593);
  not gc593 (wc593, n_1386);
  and g2254 (n_1975, n_1373, wc594);
  not gc594 (wc594, n_1374);
  and g2255 (n_1475, n_1459, wc595);
  not gc595 (wc595, n_1460);
  and g2256 (n_1976, n_1969, wc596);
  not gc596 (wc596, n_1466);
  and g2257 (n_1977, n_1453, wc597);
  not gc597 (wc597, n_1454);
  or g2258 (n_1978, wc598, n_1316);
  not gc598 (wc598, n_1315);
  or g2259 (n_1979, wc599, n_1388);
  not gc599 (wc599, n_1383);
  or g2260 (n_1980, wc600, n_1468);
  not gc600 (wc600, n_1463);
  or g2261 (n_1981, n_1308, wc601);
  not gc601 (wc601, n_1303);
  or g2262 (n_1982, n_1376, wc602);
  not gc602 (wc602, n_1371);
  or g2263 (n_1983, n_1456, wc603);
  not gc603 (wc603, n_1451);
  or g2264 (n_1984, n_1308, wc604);
  not gc604 (wc604, n_1317);
  or g2265 (n_1985, wc605, n_1304);
  not gc605 (wc605, n_1305);
  or g2266 (n_1986, n_1376, wc606);
  not gc606 (wc606, n_1389);
  or g2267 (n_1987, wc607, n_1372);
  not gc607 (wc607, n_1373);
  or g2268 (n_1988, n_1456, wc608);
  not gc608 (wc608, n_1469);
  or g2269 (n_1989, wc609, n_1452);
  not gc609 (wc609, n_1453);
  or g2270 (n_1990, n_1314, wc610);
  not gc610 (wc610, n_1309);
  or g2271 (n_1991, n_1382, wc611);
  not gc611 (wc611, n_1377);
  or g2272 (n_1992, n_1462, wc612);
  not gc612 (wc612, n_1457);
  or g2273 (n_1993, wc613, n_1310);
  not gc613 (wc613, n_1311);
  or g2274 (n_1994, wc614, n_1378);
  not gc614 (wc614, n_1379);
  or g2275 (n_1995, wc615, n_1458);
  not gc615 (wc615, n_1459);
  and g2276 (n_1996, wc616, n_1400);
  not gc616 (wc616, n_1395);
  and g2277 (n_1997, wc617, n_1480);
  not gc617 (wc617, n_1475);
  and g2278 (n_1998, n_1971, wc618);
  not gc618 (wc618, n_1329);
  or g2279 (n_1999, n_1973, wc619);
  not gc619 (wc619, n_1331);
  and g2280 (n_2000, wc620, n_1974);
  not gc620 (wc620, n_1996);
  or g2281 (n_2001, n_1413, wc621);
  not gc621 (wc621, n_1405);
  and g2282 (n_2002, wc622, n_1976);
  not gc622 (wc622, n_1997);
  or g2283 (n_2003, n_1493, wc623);
  not gc623 (wc623, n_1485);
  or g2284 (n_2004, n_1314, wc624);
  not gc624 (wc624, n_1331);
  or g2285 (n_2005, n_1382, wc625);
  not gc625 (wc625, n_1405);
  or g2286 (n_2006, n_1462, wc626);
  not gc626 (wc626, n_1485);
  or g2287 (n_2007, n_1970, wc627);
  not gc627 (wc627, n_1498);
  or g2288 (n_1297, n_1340, n_206);
  or g2289 (n_1365, n_1417, n_206);
  and g2290 (n_237, wc628, n_1297);
  not gc628 (wc628, n_1365);
  and g2291 (n_240, n_1365, wc629);
  not gc629 (wc629, n_241);
  or g2292 (n_251, wc630, wc632, wc633, wc634);
  and gc634 (wc634, n_227, n_241);
  and gc633 (wc633, n_240, n_226);
  and gc632 (wc632, n_237, n_225);
  and gc631 (wc630, wc631, n_204);
  not gc630 (wc631, n_1297);
  or g2293 (n_247, wc635, wc637, wc638, wc639);
  and gc639 (wc639, n_215, n_241);
  and gc638 (wc638, n_240, n_214);
  and gc637 (wc637, n_237, n_213);
  and gc636 (wc635, wc636, n_200);
  not gc635 (wc636, n_1297);
  or g2294 (n_248, wc640, wc642, wc643, wc644);
  and gc644 (wc644, n_218, n_241);
  and gc643 (wc643, n_240, n_217);
  and gc642 (wc642, n_237, n_216);
  and gc641 (wc640, wc641, n_201);
  not gc640 (wc641, n_1297);
  or g2295 (n_249, wc645, wc647, wc648, wc649);
  and gc649 (wc649, n_221, n_241);
  and gc648 (wc648, n_240, n_220);
  and gc647 (wc647, n_237, n_219);
  and gc646 (wc645, wc646, n_202);
  not gc645 (wc646, n_1297);
  or g2296 (n_250, wc650, wc652, wc653, wc654);
  and gc654 (wc654, n_224, n_241);
  and gc653 (wc653, n_240, n_223);
  and gc652 (wc652, n_237, n_222);
  and gc651 (wc650, wc651, n_203);
  not gc650 (wc651, n_1297);
  or g2297 (n_245, wc655, wc657, wc659, wc660);
  and gc661 (wc660, wc661, n_241);
  not gc660 (wc661, n_1764);
  and gc659 (wc659, A[2], n_240);
  and gc658 (wc657, n_237, wc658);
  not gc657 (wc658, n_1764);
  and gc656 (wc655, A[2], wc656);
  not gc655 (wc656, n_1297);
  or g2298 (n_246, wc662, wc664, wc665, wc666);
  and gc666 (wc666, n_212, n_241);
  and gc665 (wc665, n_240, n_1801);
  and gc664 (wc664, n_237, n_210);
  and gc663 (wc662, A[3], wc663);
  not gc662 (wc663, n_1297);
  or g2299 (n_1538, B[4], wc667);
  not gc667 (wc667, n_247);
  and g2300 (n_1539, B[5], wc668);
  not gc668 (wc668, n_248);
  or g2301 (n_1540, B[5], wc669);
  not gc669 (wc669, n_248);
  and g2302 (n_1545, B[6], wc670);
  not gc670 (wc670, n_249);
  or g2303 (n_1544, B[6], wc671);
  not gc671 (wc671, n_249);
  or g2304 (n_1532, B[2], wc672);
  not gc672 (wc672, n_245);
  and g2305 (n_1533, B[3], wc673);
  not gc673 (wc673, n_246);
  or g2306 (n_1534, B[3], wc674);
  not gc674 (wc674, n_246);
  and g2307 (n_1537, B[2], wc675);
  not gc675 (wc675, n_245);
  and g2308 (n_1543, B[4], wc676);
  not gc676 (wc676, n_247);
  or g2309 (n_1606, B[3], wc677);
  not gc677 (wc677, n_247);
  and g2310 (n_1607, B[4], wc678);
  not gc678 (wc678, n_248);
  or g2311 (n_1608, B[4], wc679);
  not gc679 (wc679, n_248);
  and g2312 (n_1617, B[5], wc680);
  not gc680 (wc680, n_249);
  and g2313 (n_1613, B[6], wc681);
  not gc681 (wc681, n_250);
  or g2314 (n_1612, B[5], wc682);
  not gc682 (wc682, n_249);
  or g2315 (n_2008, B[6], wc683);
  not gc683 (wc683, n_250);
  or g2316 (n_1600, B[1], wc684);
  not gc684 (wc684, n_245);
  and g2317 (n_1601, B[2], wc685);
  not gc685 (wc685, n_246);
  or g2318 (n_1602, B[2], wc686);
  not gc686 (wc686, n_246);
  and g2319 (n_1605, B[1], wc687);
  not gc687 (wc687, n_245);
  and g2320 (n_1611, B[3], wc688);
  not gc688 (wc688, n_247);
  or g2321 (n_2009, wc689, n_1823);
  not gc689 (wc689, n_251);
  or g2322 (n_1686, wc690, n_37);
  not gc690 (wc690, n_247);
  and g2323 (n_1687, wc691, n_38);
  not gc691 (wc691, n_248);
  or g2324 (n_1688, wc692, n_38);
  not gc692 (wc692, n_248);
  and g2325 (n_1697, wc693, n_39);
  not gc693 (wc693, n_249);
  and g2326 (n_1693, wc694, n_40);
  not gc694 (wc694, n_250);
  or g2327 (n_1692, wc695, n_39);
  not gc695 (wc695, n_249);
  or g2328 (n_2010, wc696, n_40);
  not gc696 (wc696, n_250);
  or g2329 (n_1680, wc697, n_1783);
  not gc697 (wc697, n_245);
  and g2330 (n_1681, wc698, n_36);
  not gc698 (wc698, n_246);
  or g2331 (n_1682, wc699, n_36);
  not gc699 (wc699, n_246);
  and g2332 (n_1685, wc700, n_1783);
  not gc700 (wc700, n_245);
  and g2333 (n_1691, wc701, n_37);
  not gc701 (wc701, n_247);
  and g2334 (n_2011, wc702, n_1823);
  not gc702 (wc702, n_251);
  and g2335 (n_1552, n_1540, wc703);
  not gc703 (wc703, n_1541);
  and g2336 (n_2012, n_1544, wc704);
  not gc704 (wc704, n_250);
  and g2337 (n_2013, n_1534, wc705);
  not gc705 (wc705, n_1535);
  or g2338 (n_2014, n_1545, wc706);
  not gc706 (wc706, n_1555);
  and g2339 (n_1624, n_1608, wc707);
  not gc707 (wc707, n_1609);
  and g2340 (n_2015, n_2008, wc708);
  not gc708 (wc708, n_1615);
  and g2341 (n_2016, n_1602, wc709);
  not gc709 (wc709, n_1603);
  and g2342 (n_1704, n_1688, wc710);
  not gc710 (wc710, n_1689);
  and g2343 (n_2017, n_2010, wc711);
  not gc711 (wc711, n_1695);
  and g2344 (n_2018, n_1682, wc712);
  not gc712 (wc712, n_1683);
  or g2345 (n_2019, n_1537, wc713);
  not gc713 (wc713, n_1546);
  or g2346 (n_2020, n_1537, wc714);
  not gc714 (wc714, n_1532);
  or g2347 (n_2021, wc715, n_1533);
  not gc715 (wc715, n_1534);
  or g2348 (n_2022, n_1543, wc716);
  not gc716 (wc716, n_1538);
  or g2349 (n_2023, wc717, n_1539);
  not gc717 (wc717, n_1540);
  or g2350 (n_2024, wc718, n_1545);
  not gc718 (wc718, n_1544);
  or g2351 (n_2025, n_1605, wc719);
  not gc719 (wc719, n_1618);
  or g2352 (n_2026, n_1605, wc720);
  not gc720 (wc720, n_1600);
  or g2353 (n_2027, wc721, n_1601);
  not gc721 (wc721, n_1602);
  or g2354 (n_2028, n_1611, wc722);
  not gc722 (wc722, n_1606);
  or g2355 (n_2029, wc723, n_1607);
  not gc723 (wc723, n_1608);
  or g2356 (n_2030, wc724, n_1617);
  not gc724 (wc724, n_1612);
  or g2357 (n_2031, n_1685, wc725);
  not gc725 (wc725, n_1698);
  or g2358 (n_2032, n_1685, wc726);
  not gc726 (wc726, n_1680);
  or g2359 (n_2033, wc727, n_1681);
  not gc727 (wc727, n_1682);
  or g2360 (n_2034, n_1691, wc728);
  not gc728 (wc728, n_1686);
  or g2361 (n_2035, wc729, n_1687);
  not gc729 (wc729, n_1688);
  or g2362 (n_2036, wc730, n_1697);
  not gc730 (wc730, n_1692);
  and g2363 (n_2037, wc731, n_1629);
  not gc731 (wc731, n_1624);
  and g2364 (n_2038, wc732, n_1709);
  not gc732 (wc732, n_1704);
  and g2365 (n_2039, n_2012, wc733);
  not gc733 (wc733, n_1558);
  or g2366 (n_2040, n_2014, wc734);
  not gc734 (wc734, n_1560);
  and g2367 (n_2041, wc735, n_2015);
  not gc735 (wc735, n_2037);
  or g2368 (n_2042, n_1642, wc736);
  not gc736 (wc736, n_1634);
  and g2369 (n_2043, wc737, n_2017);
  not gc737 (wc737, n_2038);
  or g2370 (n_2044, n_1722, wc738);
  not gc738 (wc738, n_1714);
  or g2371 (n_2045, n_1543, wc739);
  not gc739 (wc739, n_1560);
  or g2372 (n_2046, n_1611, wc740);
  not gc740 (wc740, n_1634);
  or g2373 (n_2047, n_1691, wc741);
  not gc741 (wc741, n_1714);
  or g2374 (n_2048, n_2011, wc742);
  not gc742 (wc742, n_1727);
  or g2375 (n_1526, n_1569, n_251);
  or g2376 (n_1594, n_1646, n_251);
  and g2377 (n_282, wc743, n_1526);
  not gc743 (wc743, n_1594);
  and g2378 (n_285, n_1594, wc744);
  not gc744 (wc744, n_286);
  or g2379 (REMAINDER[6], wc745, wc747, wc748, wc749);
  and gc749 (wc749, n_272, n_286);
  and gc748 (wc748, n_285, n_271);
  and gc747 (wc747, n_282, n_270);
  and gc746 (wc745, wc746, n_249);
  not gc745 (wc746, n_1526);
  or g2380 (REMAINDER[5], wc750, wc752, wc753, wc754);
  and gc754 (wc754, n_269, n_286);
  and gc753 (wc753, n_285, n_268);
  and gc752 (wc752, n_282, n_267);
  and gc751 (wc750, wc751, n_248);
  not gc750 (wc751, n_1526);
  or g2381 (REMAINDER[4], wc755, wc757, wc758, wc759);
  and gc759 (wc759, n_266, n_286);
  and gc758 (wc758, n_285, n_265);
  and gc757 (wc757, n_282, n_264);
  and gc756 (wc755, wc756, n_247);
  not gc755 (wc756, n_1526);
  or g2382 (REMAINDER[3], wc760, wc762, wc763, wc764);
  and gc764 (wc764, n_263, n_286);
  and gc763 (wc763, n_285, n_262);
  and gc762 (wc762, n_282, n_261);
  and gc761 (wc760, wc761, n_246);
  not gc760 (wc761, n_1526);
  or g2383 (REMAINDER[2], wc765, wc767, wc768, wc769);
  and gc769 (wc769, n_260, n_286);
  and gc768 (wc768, n_285, n_259);
  and gc767 (wc767, n_282, n_258);
  and gc766 (wc765, wc766, n_245);
  not gc765 (wc766, n_1526);
  or g2384 (REMAINDER[1], wc770, wc772, wc773, wc774);
  and gc774 (wc774, n_257, n_286);
  and gc773 (wc773, n_285, n_1804);
  and gc772 (wc772, n_282, n_255);
  and gc771 (wc770, A[1], wc771);
  not gc770 (wc771, n_1526);
  or g2385 (REMAINDER[0], wc775, wc777, wc779, wc780);
  and gc781 (wc780, wc781, n_286);
  not gc780 (wc781, n_1766);
  and gc779 (wc779, A[0], n_285);
  and gc778 (wc777, n_282, wc778);
  not gc777 (wc778, n_1766);
  and gc776 (wc775, A[0], wc776);
  not gc775 (wc776, n_1526);
endmodule

module remainder_unsigned_268_GENERIC(A, B, REMAINDER);
  input [14:0] A;
  input [6:0] B;
  output [14:0] REMAINDER;
  wire [14:0] A;
  wire [6:0] B;
  wire [14:0] REMAINDER;
  remainder_unsigned_268_GENERIC_REAL g1(.A (A), .B (B), .REMAINDER
       (REMAINDER));
endmodule

